* First line

.INCLUDE "cmosedu_models.txt"

.MODEL NMOS NMOS
.MODEL PMOS PMOS

.GLOBAL vdd!

*.TEMP 25.0

*.OPTION INGOLD=2 ARTIST=2 PSF=2 MEASOUT=1 PARHIER=LOCAL PROBE=0 MARCH=2 ACCURACY=1 POST

.SUBCKT nmos_rvt d g s b PARAMS: w=270e-9 l=20e-9 nfin=12
.param width={nfin*200n}
.param length={50n}
.param perimeter={3*length}
.param area={1.5*length*width}

mn d g s b N_50n L={length} W={width} PD={perimeter} AD={area}
.ENDS

.SUBCKT pmos_rvt d g s b PARAMS: w=270e-9 l=20e-9 nfin=12
.param width={nfin*200n}
.param length={50n}
.param perimeter={3*length}
.param area={1.5*length*width}

mp d g s b P_50n L={length} W={width} PD={perimeter} AD={area}
.ENDS

r698 net_m1_M1_X0_Y0_G net8 50
r699 net_m1_M1_X0_Y0_S vdd! 50
r700 net_m1_M1_X0_Y0_S vdd! 50
r701 net_m1_M1_X0_Y0_S vdd! 50
r702 net_m1_M1_X0_Y0_D net8 50
r703 net_m1_M1_X0_Y0_D net8 50
r704 net_m1_M1_X0_Y0_D net8 50
r705 net_m2_M1_X0_Y0_G net8 50
r706 net_m2_M1_X0_Y0_S vdd! 50
r707 net_m2_M1_X0_Y0_S vdd! 50
r708 net_m2_M1_X0_Y0_S vdd! 50
r709 net_m2_M1_X0_Y0_D vout 50
r710 net_m2_M1_X0_Y0_D vout 50
r711 net_m2_M1_X0_Y0_D vout 50
r712 net_m5_m4_M1_X0_Y0_G id 50
r713 net_m5_m4_M1_X0_Y0_S 0 50
r714 net_m5_m4_M1_X0_Y0_S 0 50
r715 net_m5_m4_M1_X0_Y0_S 0 50
r716 net_m5_m4_M1_X0_Y0_D id 50
r717 net_m5_m4_M1_X0_Y0_D id 50
r718 net_m5_m4_M1_X0_Y0_D id 50
r719 net_m5_m4_M2_X1_Y0_G id 50
r720 net_m5_m4_M2_X1_Y0_S 0 50
r721 net_m5_m4_M2_X1_Y0_S 0 50
r722 net_m5_m4_M2_X1_Y0_S 0 50
r723 net_m5_m4_M2_X1_Y0_D net10 50
r724 net_m5_m4_M2_X1_Y0_D net10 50
r725 net_m5_m4_M2_X1_Y0_D net10 50
r726 net_m0_m3_M1_X0_Y0_G vinp 50
r727 net_m0_m3_M1_X0_Y0_S net10 50
r728 net_m0_m3_M1_X0_Y0_S net10 50
r729 net_m0_m3_M1_X0_Y0_S net10 50
r730 net_m0_m3_M1_X0_Y0_D net8 50
r731 net_m0_m3_M1_X0_Y0_D net8 50
r732 net_m0_m3_M1_X0_Y0_D net8 50
r733 net_m0_m3_M2_X1_Y0_G vinn 50
r734 net_m0_m3_M2_X1_Y0_S net10 50
r735 net_m0_m3_M2_X1_Y0_S net10 50
r736 net_m0_m3_M2_X1_Y0_S net10 50
r737 net_m0_m3_M2_X1_Y0_D vout 50
r738 net_m0_m3_M2_X1_Y0_D vout 50
r739 net_m0_m3_M2_X1_Y0_D vout 50

x_m1_M1_X0_Y0_0 net_m1_M1_X0_Y0_D net_m1_M1_X0_Y0_G net_m1_M1_X0_Y0_diff vdd! pmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m1_M1_X0_Y0_1 net_m1_M1_X0_Y0_diff net_m1_M1_X0_Y0_G net_m1_M1_X0_Y0_S vdd! pmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m2_M1_X0_Y0_0 net_m2_M1_X0_Y0_D net_m2_M1_X0_Y0_G net_m2_M1_X0_Y0_diff vdd! pmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m2_M1_X0_Y0_1 net_m2_M1_X0_Y0_diff net_m2_M1_X0_Y0_G net_m2_M1_X0_Y0_S vdd! pmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m5_m4_M1_X0_Y0_0 net_m5_m4_M1_X0_Y0_D net_m5_m4_M1_X0_Y0_G net_m5_m4_M1_X0_Y0_diff gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m5_m4_M1_X0_Y0_1 net_m5_m4_M1_X0_Y0_diff net_m5_m4_M1_X0_Y0_G net_m5_m4_M1_X0_Y0_S gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m5_m4_M2_X1_Y0_0 net_m5_m4_M2_X1_Y0_D net_m5_m4_M2_X1_Y0_G net_m5_m4_M2_X1_Y0_diff gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m5_m4_M2_X1_Y0_1 net_m5_m4_M2_X1_Y0_diff net_m5_m4_M2_X1_Y0_G net_m5_m4_M2_X1_Y0_S gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m0_m3_M1_X0_Y0_0 net_m0_m3_M1_X0_Y0_D net_m0_m3_M1_X0_Y0_G net_m0_m3_M1_X0_Y0_diff gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m0_m3_M1_X0_Y0_1 net_m0_m3_M1_X0_Y0_diff net_m0_m3_M1_X0_Y0_G net_m0_m3_M1_X0_Y0_S gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m0_m3_M2_X1_Y0_0 net_m0_m3_M2_X1_Y0_D net_m0_m3_M2_X1_Y0_G net_m0_m3_M2_X1_Y0_diff gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m0_m3_M2_X1_Y0_1 net_m0_m3_M2_X1_Y0_diff net_m0_m3_M2_X1_Y0_G net_m0_m3_M2_X1_Y0_S gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12

**testbench
v2 vinp 0 DC 675e-3 AC .5 180 SIN(675e-3 .002 1k 0 0 180)
v1 vinn 0 DC 675e-3 AC .5     SIN(675e-3 .002 1k 0 0   0)
v0 vdd! 0 1.0
i5 vdd! id 40e-6
cload vout 0 350e-15

*.OP

*.PRINT DC v(vout) v(id) v(vinp) v(vinn) id(x_m5_m4_M2_X1_Y0_0:mn) id(x_m5_m4_M2_X1_Y0_1:mn) id(x_m5_m4_M1_X0_Y0_0:mn) id(x_m5_m4_M1_X0_Y0_1:mn)

.AC DEC 100 1.0 1e11
.PRINT AC vdb(vout) vm(vout)

*.tran 10n 5m
*.PRINT TRAN v(vout) v(vinp) v(vinn) v(id) v(net10) v(net8)
*.OPTIONS OUTPUT INITIAL_INTERVAL=1u
*.OPTIONS TIMEINT RELTOL=1e-4 ABSTOL=1e-8

*.MEASURE TRAN vout_max MAX v(vout)
*.MEASURE TRAN vout_min MIN v(vout)
*.MEASURE TRAN vout_pp  PP  v(vout)

.END

*
* Short channel models from CMOS Circuit Design, Layout, and Simulation,
* 50nm BSIM4 models VDD=1V, see CMOSedu.com
*
.model  N_50n  nmos  level = 54
+binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 0          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0          
+tnom    = 27           toxe    = 1.4e-009     toxp    = 7e-010       toxm    = 1.4e-009   
+epsrox  = 3.9          wint    = 5e-009       lint    = 1.2e-008   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 1.4e-009   
+vth0    = 0.22         k1      = 0.35         k2      = 0.05         k3      = 0          
+k3b     = 0            w0      = 2.5e-006     dvt0    = 2.8          dvt1    = 0.52       
+dvt2    = -0.032       dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 2            minv    = 0.05         voffl   = 0            dvtp0   = 1e-007     
+dvtp1   = 0.05         lpe0    = 5.75e-008    lpeb    = 2.3e-010     xj      = 2e-008     
+ngate   = 5e+020       ndep    = 2.8e+018     nsd     = 1e+020       phin    = 0          
+cdsc    = 0.0002       cdscb   = 0            cdscd   = 0            cit     = 0          
+voff    = -0.15        nfactor = 1.2          eta0    = 0.15         etab    = 0          
+vfb     = -0.55        u0      = 0.032        ua      = 1.6e-010     ub      = 1.1e-017   
+uc      = -3e-011      vsat    = 1.1e+005     a0      = 2            ags     = 1e-020     
+a1      = 0            a2      = 1            b0      = -1e-020      b1      = 0          
+keta    = 0.04         dwg     = 0            dwb     = 0            pclm    = 0.18       
+pdiblc1 = 0.028        pdiblc2 = 0.022        pdiblcb = -0.005       drout   = 0.45       
+pvag    = 1e-020       delta   = 0.01         pscbe1  = 8.14e+008    pscbe2  = 1e-007     
+fprout  = 0.2          pdits   = 0.2          pditsd  = 0.23         pditsl  = 2.3e+006   
+rsh     = 3            rdsw    = 150          rsw     = 150          rdw     = 150        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 0          
+prwb    = 6.8e-011     wr      = 1            alpha0  = 0.074        alpha1  = 0.005      
+beta0   = 30           agidl   = 0.0002       bgidl   = 2.1e+009     cgidl   = 0.0002     
+egidl   = 0.8          
+aigbacc = 0.012        bigbacc = 0.0028       cigbacc = 0.002
+nigbacc = 1            aigbinv = 0.014        bigbinv = 0.004        cigbinv = 0.004
+eigbinv = 1.1          nigbinv = 3            aigc    = 0.017        bigc    = 0.0028
+cigc    = 0.002        aigsd   = 0.017        bigsd   = 0.0028       cigsd   = 0.002
+nigc    = 1            poxedge = 1            pigcd   = 1            ntox    = 1
+xrcrg1  = 12           xrcrg2  = 5          
+cgso    = 6.238e-010   cgdo    = 6.238e-010   cgbo    = 2.56e-011    cgdl    = 2.495e-10     
+cgsl    = 2.495e-10    ckappas = 0.02         ckappad = 0.02         acde    = 1          
+moin    = 15           noff    = 0.9          voffcv  = 0.02       
+kt1     = -0.21        kt1l    = 0.0           kt2     = -0.042        ute     = -1.5
+ua1     = 1e-009       ub1     = -3.5e-019     uc1     = 0             prt     = 0
+at      = 53000
+fnoimod = 1            tnoimod = 0          
+jss     = 0.0001       jsws    = 1e-011       jswgs   = 1e-010       njs     = 1          
+ijthsfwd= 0.01         ijthsrev= 0.001        bvs     = 10           xjbvs   = 1          
+jsd     = 0.0001       jswd    = 1e-011       jswgd   = 1e-010       njd     = 1          
+ijthdfwd= 0.01         ijthdrev= 0.001        bvd     = 10           xjbvd   = 1          
+pbs     = 1            cjs     = 0.0005       mjs     = 0.5          pbsws   = 1          
+cjsws   = 5e-010       mjsws   = 0.33         pbswgs  = 1            cjswgs  = 5e-010     
+mjswgs  = 0.33         pbd     = 1            cjd     = 0.0005       mjd     = 0.5        
+pbswd   = 1            cjswd   = 5e-010       mjswd   = 0.33         pbswgd  = 1          
+cjswgd  = 5e-010       mjswgd  = 0.33         tpb     = 0.005        tcj     = 0.001      
+tpbsw   = 0.005        tcjsw   = 0.001        tpbswg  = 0.005        tcjswg  = 0.001      
+xtis    = 3            xtid    = 3          
+dmcg    = 0e-006       dmci    = 0e-006       dmdg    = 0e-006       dmcgt   = 0e-007     
+dwj     = 0e-008     	xgw     = 0e-007       xgl     = 0e-008     
+rshg    = 0.4          gbmin   = 1e-010       rbpb    = 5            rbpd    = 15         
+rbps    = 15           rbdb    = 15           rbsb    = 15           ngcon   = 1
*
.model  P_50n  pmos  level = 54
+binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 0          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0          
+tnom    = 27           toxe    = 1.4e-009     toxp    = 7e-010       toxm    = 1.4e-009   
+epsrox  = 3.9          wint    = 5e-009       lint    = 1.2e-008   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 1.4e-009   
+vth0    = -0.22        k1      = 0.39         k2      = 0.05         k3      = 0          
+k3b     = 0            w0      = 2.5e-006     dvt0    = 3.9          dvt1    = 0.635        
+dvt2    = -0.032       dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 0.7          minv    = 0.05         voffl   = 0            dvtp0   = 0.5e-008     
+dvtp1   = 0.05         lpe0    = 5.75e-008    lpeb    = 2.3e-010     xj      = 2e-008     
+ngate   = 5e+020       ndep    = 2.8e+018     nsd     = 1e+020       phin    = 0          
+cdsc    = 0.000258     cdscb   = 0            cdscd   = 6.1e-008     cit     = 0          
+voff    = -0.15        nfactor = 2            eta0    = 0.15         etab    = 0          
+vfb     = 0.55         u0      = 0.0095       ua      = 1.6e-009     ub      = 8e-018     
+uc      = 4.6e-013     vsat    = 90000        a0      = 1.2          ags     = 1e-020     
+a1      = 0            a2      = 1            b0      = -1e-020      b1      = 0          
+keta    = -0.047       dwg     = 0            dwb     = 0            pclm    = 0.55       
+pdiblc1 = 0.03         pdiblc2 = 0.0055       pdiblcb = 3.4e-008     drout   = 0.56       
+pvag    = 1e-020       delta   = 0.014        pscbe1  = 8.14e+008    pscbe2  = 9.58e-007  
+fprout  = 0.2          pdits   = 0.2          pditsd  = 0.23         pditsl  = 2.3e+006   
+rsh     = 3            rdsw    = 250          rsw     = 160          rdw     = 160        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 3.22e-008  
+prwb    = 6.8e-011     wr      = 1            alpha0  = 0.074        alpha1  = 0.005      
+beta0   = 30           agidl   = 0.0002       bgidl   = 2.1e+009     cgidl   = 0.0002     
+egidl   = 0.8          
+aigbacc = 0.012        bigbacc = 0.0028       cigbacc = 0.002
+nigbacc = 1            aigbinv = 0.014        bigbinv = 0.004        cigbinv = 0.004
+eigbinv = 1.1          nigbinv = 3            aigc    = 0.69         bigc    = 0.0012
+cigc    = 0.0008       aigsd   = 0.0087       bigsd   = 0.0012       cigsd   = 0.0008
+nigc    = 1            poxedge = 1            pigcd   = 1            ntox    = 1
+xrcrg1  = 12           xrcrg2  = 5          
+cgso    = 7.43e-010    cgdo    = 7.43e-010    cgbo    = 2.56e-011    cgdl    = 1e-014     
+cgsl    = 1e-014       ckappas = 0.5          ckappad = 0.5          acde    = 1          
+moin    = 15           noff    = 0.9          voffcv  = 0.02       
+kt1     = -0.19        kt1l    = 0            kt2     = -0.052        ute     = -1.5
+ua1     = -1e-009      ub1     = 2e-018       uc1     = 0             prt     = 0
+at      = 33000
+fnoimod = 1            tnoimod = 0          
+jss     = 0.0001       jsws    = 1e-011       jswgs   = 1e-010       njs     = 1          
+ijthsfwd= 0.01         ijthsrev= 0.001        bvs     = 10           xjbvs   = 1          
+jsd     = 0.0001       jswd    = 1e-011       jswgd   = 1e-010       njd     = 1          
+ijthdfwd= 0.01         ijthdrev= 0.001        bvd     = 10           xjbvd   = 1          
+pbs     = 1            cjs     = 0.0005       mjs     = 0.5          pbsws   = 1          
+cjsws   = 5e-010       mjsws   = 0.33         pbswgs  = 1            cjswgs  = 5e-010     
+mjswgs  = 0.33         pbd     = 1            cjd     = 0.0005       mjd     = 0.5        
+pbswd   = 1            cjswd   = 5e-010       mjswd   = 0.33         pbswgd  = 1          
+cjswgd  = 5e-010       mjswgd  = 0.33         tpb     = 0.005        tcj     = 0.001      
+tpbsw   = 0.005        tcjsw   = 0.001        tpbswg  = 0.005        tcjswg  = 0.001      
+xtis    = 3            xtid    = 3          
+dmcg    = 0e-006       dmci    = 0e-006       dmdg    = 0e-006       dmcgt   = 0e-007     
+dwj     = 0e-008     	xgw     = 0e-007       xgl     = 0e-008     
+rshg    = 0.4          gbmin   = 1e-010       rbpb    = 5            rbpd    = 15         
+rbps    = 15           rbdb    = 15           rbsb    = 15           ngcon   = 1   


.MODEL NMOS NMOS
.MODEL PMOS PMOS

.GLOBAL vdd!

*.TEMP 25.0

*.OPTION INGOLD=2 ARTIST=2 PSF=2 MEASOUT=1 PARHIER=LOCAL PROBE=0 MARCH=2 ACCURACY=1 POST

.SUBCKT nmos_rvt d g s b PARAMS: w=270e-9 l=20e-9 nfin=12
.param width={nfin*200n}
.param length={50n}
.param perimeter={3*length}
.param area={1.5*length*width}

mn d g s b N_50n L={length} W={width} PD={perimeter} AD={area}
.ENDS

.SUBCKT pmos_rvt d g s b PARAMS: w=270e-9 l=20e-9 nfin=12
.param width={nfin*200n}
.param length={50n}
.param perimeter={3*length}
.param area={1.5*length*width}

mp d g s b P_50n L={length} W={width} PD={perimeter} AD={area}
.ENDS

r0 net8_M1_3840_132 net8_M1_3840_168 3.5999999999999996
c0 net8_M1_3840_132 0 0.0036f
c1 net8_M1_3840_168 0 0.0036f
r1 net8_M1_3840_168 net8_M1_3840_248 8.0
c2 net8_M1_3840_168 0 0.008f
c3 net8_M1_3840_248 0 0.008f
r2 net8_M1_3840_248 net8_M1_3840_252 0.4
c4 net8_M1_3840_248 0 0.0004f
c5 net8_M1_3840_252 0 0.0004f
r3 net8_M1_3840_252 net8_M1_3840_332 8.0
c6 net8_M1_3840_252 0 0.008f
c7 net8_M1_3840_332 0 0.008f
r4 net8_M1_3840_332 net8_M1_3840_412 8.0
c8 net8_M1_3840_332 0 0.008f
c9 net8_M1_3840_412 0 0.008f
r5 net8_M1_3840_412 net8_M1_3840_420 0.8
c10 net8_M1_3840_412 0 0.0008f
c11 net8_M1_3840_420 0 0.0008f
r6 net8_M1_3840_420 net8_M1_3840_500 8.0
c12 net8_M1_3840_420 0 0.008f
c13 net8_M1_3840_500 0 0.008f
r7 net8_M1_3840_500 net8_M1_3840_580 8.0
c14 net8_M1_3840_500 0 0.008f
c15 net8_M1_3840_580 0 0.008f
r8 net8_M1_3840_580 net8_M1_3840_660 8.0
c16 net8_M1_3840_580 0 0.008f
c17 net8_M1_3840_660 0 0.008f
r9 net8_M1_3840_660 net8_M1_3840_740 8.0
c18 net8_M1_3840_660 0 0.008f
c19 net8_M1_3840_740 0 0.008f
r10 net8_M1_3840_740 net8_M1_3840_792 5.2
c20 net8_M1_3840_740 0 0.0052f
c21 net8_M1_3840_792 0 0.0052f
r11 vdd_M1_3920_132 vdd_M1_3920_168 3.5999999999999996
c22 vdd_M1_3920_132 0 0.0036f
c23 vdd_M1_3920_168 0 0.0036f
r12 vdd_M1_3920_168 vdd_M1_3920_248 8.0
c24 vdd_M1_3920_168 0 0.008f
c25 vdd_M1_3920_248 0 0.008f
r13 vdd_M1_3920_248 vdd_M1_3920_328 8.0
c26 vdd_M1_3920_248 0 0.008f
c27 vdd_M1_3920_328 0 0.008f
r14 vdd_M1_3920_328 vdd_M1_3920_336 0.8
c28 vdd_M1_3920_328 0 0.0008f
c29 vdd_M1_3920_336 0 0.0008f
r15 vdd_M1_3920_336 vdd_M1_3920_416 8.0
c30 vdd_M1_3920_336 0 0.008f
c31 vdd_M1_3920_416 0 0.008f
r16 vdd_M1_3920_416 vdd_M1_3920_462 4.6
c32 vdd_M1_3920_416 0 0.0046f
c33 vdd_M1_3920_462 0 0.0046f
r17 vdd_M1_3920_462 vdd_M1_3920_542 8.0
c34 vdd_M1_3920_462 0 0.008f
c35 vdd_M1_3920_542 0 0.008f
r18 vdd_M1_3920_542 vdd_M1_3920_588 4.6
c36 vdd_M1_3920_542 0 0.0046f
c37 vdd_M1_3920_588 0 0.0046f
r19 vdd_M1_3920_588 vdd_M1_3920_668 8.0
c38 vdd_M1_3920_588 0 0.008f
c39 vdd_M1_3920_668 0 0.008f
r20 vdd_M1_3920_668 vdd_M1_3920_748 8.0
c40 vdd_M1_3920_668 0 0.008f
c41 vdd_M1_3920_748 0 0.008f
r21 vdd_M1_3920_748 vdd_M1_3920_792 4.3999999999999995
c42 vdd_M1_3920_748 0 0.0044f
c43 vdd_M1_3920_792 0 0.0044f
r22 net8_M1_3760_132 net8_M1_3760_212 8.0
c44 net8_M1_3760_132 0 0.008f
c45 net8_M1_3760_212 0 0.008f
r23 net8_M1_3760_212 net8_M1_3760_252 4.0
c46 net8_M1_3760_212 0 0.004f
c47 net8_M1_3760_252 0 0.004f
r24 net8_M1_3760_252 net8_M1_3760_332 8.0
c48 net8_M1_3760_252 0 0.008f
c49 net8_M1_3760_332 0 0.008f
r25 net8_M1_3760_332 net8_M1_3760_336 0.4
c50 net8_M1_3760_332 0 0.0004f
c51 net8_M1_3760_336 0 0.0004f
r26 net8_M1_3760_336 net8_M1_3760_416 8.0
c52 net8_M1_3760_336 0 0.008f
c53 net8_M1_3760_416 0 0.008f
r27 net8_M1_3760_416 net8_M1_3760_420 0.4
c54 net8_M1_3760_416 0 0.0004f
c55 net8_M1_3760_420 0 0.0004f
r28 net8_M1_3760_420 net8_M1_3760_462 4.2
c56 net8_M1_3760_420 0 0.004200000000000001f
c57 net8_M1_3760_462 0 0.004200000000000001f
r29 net8_M1_3760_462 net8_M1_3760_542 8.0
c58 net8_M1_3760_462 0 0.008f
c59 net8_M1_3760_542 0 0.008f
r30 net8_M1_3760_542 net8_M1_3760_588 4.6
c60 net8_M1_3760_542 0 0.0046f
c61 net8_M1_3760_588 0 0.0046f
r31 net8_M1_3760_588 net8_M1_3760_668 8.0
c62 net8_M1_3760_588 0 0.008f
c63 net8_M1_3760_668 0 0.008f
r32 net8_M1_3760_668 net8_M1_3760_748 8.0
c64 net8_M1_3760_668 0 0.008f
c65 net8_M1_3760_748 0 0.008f
r33 net8_M1_3760_748 net8_M1_3760_792 4.3999999999999995
c66 net8_M1_3760_748 0 0.0044f
c67 net8_M1_3760_792 0 0.0044f
r34 net8_M1_3120_132 net8_M1_3120_168 3.5999999999999996
c68 net8_M1_3120_132 0 0.0036f
c69 net8_M1_3120_168 0 0.0036f
r35 net8_M1_3120_168 net8_M1_3120_248 8.0
c70 net8_M1_3120_168 0 0.008f
c71 net8_M1_3120_248 0 0.008f
r36 net8_M1_3120_248 net8_M1_3120_328 8.0
c72 net8_M1_3120_248 0 0.008f
c73 net8_M1_3120_328 0 0.008f
r37 net8_M1_3120_328 net8_M1_3120_336 0.8
c74 net8_M1_3120_328 0 0.0008f
c75 net8_M1_3120_336 0 0.0008f
r38 net8_M1_3120_336 net8_M1_3120_416 8.0
c76 net8_M1_3120_336 0 0.008f
c77 net8_M1_3120_416 0 0.008f
r39 net8_M1_3120_416 net8_M1_3120_496 8.0
c78 net8_M1_3120_416 0 0.008f
c79 net8_M1_3120_496 0 0.008f
r40 net8_M1_3120_496 net8_M1_3120_576 8.0
c80 net8_M1_3120_496 0 0.008f
c81 net8_M1_3120_576 0 0.008f
r41 net8_M1_3120_576 net8_M1_3120_588 1.2
c82 net8_M1_3120_576 0 0.0012000000000000001f
c83 net8_M1_3120_588 0 0.0012000000000000001f
r42 net8_M1_3120_588 net8_M1_3120_668 8.0
c84 net8_M1_3120_588 0 0.008f
c85 net8_M1_3120_668 0 0.008f
r43 net8_M1_3120_668 net8_M1_3120_748 8.0
c86 net8_M1_3120_668 0 0.008f
c87 net8_M1_3120_748 0 0.008f
r44 net8_M1_3120_748 net8_M1_3120_792 4.3999999999999995
c88 net8_M1_3120_748 0 0.0044f
c89 net8_M1_3120_792 0 0.0044f
r45 vdd_M1_3200_132 vdd_M1_3200_168 3.5999999999999996
c90 vdd_M1_3200_132 0 0.0036f
c91 vdd_M1_3200_168 0 0.0036f
r46 vdd_M1_3200_168 vdd_M1_3200_248 8.0
c92 vdd_M1_3200_168 0 0.008f
c93 vdd_M1_3200_248 0 0.008f
r47 vdd_M1_3200_248 vdd_M1_3200_328 8.0
c94 vdd_M1_3200_248 0 0.008f
c95 vdd_M1_3200_328 0 0.008f
r48 vdd_M1_3200_328 vdd_M1_3200_336 0.8
c96 vdd_M1_3200_328 0 0.0008f
c97 vdd_M1_3200_336 0 0.0008f
r49 vdd_M1_3200_336 vdd_M1_3200_416 8.0
c98 vdd_M1_3200_336 0 0.008f
c99 vdd_M1_3200_416 0 0.008f
r50 vdd_M1_3200_416 vdd_M1_3200_420 0.4
c100 vdd_M1_3200_416 0 0.0004f
c101 vdd_M1_3200_420 0 0.0004f
r51 vdd_M1_3200_420 vdd_M1_3200_462 4.2
c102 vdd_M1_3200_420 0 0.004200000000000001f
c103 vdd_M1_3200_462 0 0.004200000000000001f
r52 vdd_M1_3200_462 vdd_M1_3200_542 8.0
c104 vdd_M1_3200_462 0 0.008f
c105 vdd_M1_3200_542 0 0.008f
r53 vdd_M1_3200_542 vdd_M1_3200_588 4.6
c106 vdd_M1_3200_542 0 0.0046f
c107 vdd_M1_3200_588 0 0.0046f
r54 vdd_M1_3200_588 vdd_M1_3200_668 8.0
c108 vdd_M1_3200_588 0 0.008f
c109 vdd_M1_3200_668 0 0.008f
r55 vdd_M1_3200_668 vdd_M1_3200_748 8.0
c110 vdd_M1_3200_668 0 0.008f
c111 vdd_M1_3200_748 0 0.008f
r56 vdd_M1_3200_748 vdd_M1_3200_792 4.3999999999999995
c112 vdd_M1_3200_748 0 0.0044f
c113 vdd_M1_3200_792 0 0.0044f
r57 vout_M1_3040_132 vout_M1_3040_212 8.0
c114 vout_M1_3040_132 0 0.008f
c115 vout_M1_3040_212 0 0.008f
r58 vout_M1_3040_212 vout_M1_3040_252 4.0
c116 vout_M1_3040_212 0 0.004f
c117 vout_M1_3040_252 0 0.004f
r59 vout_M1_3040_252 vout_M1_3040_332 8.0
c118 vout_M1_3040_252 0 0.008f
c119 vout_M1_3040_332 0 0.008f
r60 vout_M1_3040_332 vout_M1_3040_336 0.4
c120 vout_M1_3040_332 0 0.0004f
c121 vout_M1_3040_336 0 0.0004f
r61 vout_M1_3040_336 vout_M1_3040_416 8.0
c122 vout_M1_3040_336 0 0.008f
c123 vout_M1_3040_416 0 0.008f
r62 vout_M1_3040_416 vout_M1_3040_462 4.6
c124 vout_M1_3040_416 0 0.0046f
c125 vout_M1_3040_462 0 0.0046f
r63 vout_M1_3040_462 vout_M1_3040_504 4.2
c126 vout_M1_3040_462 0 0.004200000000000001f
c127 vout_M1_3040_504 0 0.004200000000000001f
r64 vout_M1_3040_504 vout_M1_3040_584 8.0
c128 vout_M1_3040_504 0 0.008f
c129 vout_M1_3040_584 0 0.008f
r65 vout_M1_3040_584 vout_M1_3040_588 0.4
c130 vout_M1_3040_584 0 0.0004f
c131 vout_M1_3040_588 0 0.0004f
r66 vout_M1_3040_588 vout_M1_3040_668 8.0
c132 vout_M1_3040_588 0 0.008f
c133 vout_M1_3040_668 0 0.008f
r67 vout_M1_3040_668 vout_M1_3040_748 8.0
c134 vout_M1_3040_668 0 0.008f
c135 vout_M1_3040_748 0 0.008f
r68 vout_M1_3040_748 vout_M1_3040_792 4.3999999999999995
c136 vout_M1_3040_748 0 0.0044f
c137 vout_M1_3040_792 0 0.0044f
r69 id_M1_400_132 id_M1_400_168 3.5999999999999996
c138 id_M1_400_132 0 0.0036f
c139 id_M1_400_168 0 0.0036f
r70 id_M1_400_168 id_M1_400_248 8.0
c140 id_M1_400_168 0 0.008f
c141 id_M1_400_248 0 0.008f
r71 id_M1_400_248 id_M1_400_252 0.4
c142 id_M1_400_248 0 0.0004f
c143 id_M1_400_252 0 0.0004f
r72 id_M1_400_252 id_M1_400_332 8.0
c144 id_M1_400_252 0 0.008f
c145 id_M1_400_332 0 0.008f
r73 id_M1_400_332 id_M1_400_412 8.0
c146 id_M1_400_332 0 0.008f
c147 id_M1_400_412 0 0.008f
r74 id_M1_400_412 id_M1_400_492 8.0
c148 id_M1_400_412 0 0.008f
c149 id_M1_400_492 0 0.008f
r75 id_M1_400_492 id_M1_400_504 1.2
c150 id_M1_400_492 0 0.0012000000000000001f
c151 id_M1_400_504 0 0.0012000000000000001f
r76 id_M1_400_504 id_M1_400_584 8.0
c152 id_M1_400_504 0 0.008f
c153 id_M1_400_584 0 0.008f
r77 id_M1_400_584 id_M1_400_664 8.0
c154 id_M1_400_584 0 0.008f
c155 id_M1_400_664 0 0.008f
r78 id_M1_400_664 id_M1_400_744 8.0
c156 id_M1_400_664 0 0.008f
c157 id_M1_400_744 0 0.008f
r79 id_M1_400_744 id_M1_400_792 4.8
c158 id_M1_400_744 0 0.0048000000000000004f
c159 id_M1_400_792 0 0.0048000000000000004f
r80 vss_M1_320_132 vss_M1_320_168 3.5999999999999996
c160 vss_M1_320_132 0 0.0036f
c161 vss_M1_320_168 0 0.0036f
r81 vss_M1_320_168 vss_M1_320_248 8.0
c162 vss_M1_320_168 0 0.008f
c163 vss_M1_320_248 0 0.008f
r82 vss_M1_320_248 vss_M1_320_328 8.0
c164 vss_M1_320_248 0 0.008f
c165 vss_M1_320_328 0 0.008f
r83 vss_M1_320_328 vss_M1_320_336 0.8
c166 vss_M1_320_328 0 0.0008f
c167 vss_M1_320_336 0 0.0008f
r84 vss_M1_320_336 vss_M1_320_416 8.0
c168 vss_M1_320_336 0 0.008f
c169 vss_M1_320_416 0 0.008f
r85 vss_M1_320_416 vss_M1_320_420 0.4
c170 vss_M1_320_416 0 0.0004f
c171 vss_M1_320_420 0 0.0004f
r86 vss_M1_320_420 vss_M1_320_462 4.2
c172 vss_M1_320_420 0 0.004200000000000001f
c173 vss_M1_320_462 0 0.004200000000000001f
r87 vss_M1_320_462 vss_M1_320_542 8.0
c174 vss_M1_320_462 0 0.008f
c175 vss_M1_320_542 0 0.008f
r88 vss_M1_320_542 vss_M1_320_588 4.6
c176 vss_M1_320_542 0 0.0046f
c177 vss_M1_320_588 0 0.0046f
r89 vss_M1_320_588 vss_M1_320_668 8.0
c178 vss_M1_320_588 0 0.008f
c179 vss_M1_320_668 0 0.008f
r90 vss_M1_320_668 vss_M1_320_748 8.0
c180 vss_M1_320_668 0 0.008f
c181 vss_M1_320_748 0 0.008f
r91 vss_M1_320_748 vss_M1_320_792 4.3999999999999995
c182 vss_M1_320_748 0 0.0044f
c183 vss_M1_320_792 0 0.0044f
r92 id_M1_480_132 id_M1_480_212 8.0
c184 id_M1_480_132 0 0.008f
c185 id_M1_480_212 0 0.008f
r93 id_M1_480_212 id_M1_480_252 4.0
c186 id_M1_480_212 0 0.004f
c187 id_M1_480_252 0 0.004f
r94 id_M1_480_252 id_M1_480_332 8.0
c188 id_M1_480_252 0 0.008f
c189 id_M1_480_332 0 0.008f
r95 id_M1_480_332 id_M1_480_336 0.4
c190 id_M1_480_332 0 0.0004f
c191 id_M1_480_336 0 0.0004f
r96 id_M1_480_336 id_M1_480_416 8.0
c192 id_M1_480_336 0 0.008f
c193 id_M1_480_416 0 0.008f
r97 id_M1_480_416 id_M1_480_462 4.6
c194 id_M1_480_416 0 0.0046f
c195 id_M1_480_462 0 0.0046f
r98 id_M1_480_462 id_M1_480_504 4.2
c196 id_M1_480_462 0 0.004200000000000001f
c197 id_M1_480_504 0 0.004200000000000001f
r99 id_M1_480_504 id_M1_480_584 8.0
c198 id_M1_480_504 0 0.008f
c199 id_M1_480_584 0 0.008f
r100 id_M1_480_584 id_M1_480_588 0.4
c200 id_M1_480_584 0 0.0004f
c201 id_M1_480_588 0 0.0004f
r101 id_M1_480_588 id_M1_480_668 8.0
c202 id_M1_480_588 0 0.008f
c203 id_M1_480_668 0 0.008f
r102 id_M1_480_668 id_M1_480_748 8.0
c204 id_M1_480_668 0 0.008f
c205 id_M1_480_748 0 0.008f
r103 id_M1_480_748 id_M1_480_792 4.3999999999999995
c206 id_M1_480_748 0 0.0044f
c207 id_M1_480_792 0 0.0044f
r104 id_M1_1040_132 id_M1_1040_168 3.5999999999999996
c208 id_M1_1040_132 0 0.0036f
c209 id_M1_1040_168 0 0.0036f
r105 id_M1_1040_168 id_M1_1040_248 8.0
c210 id_M1_1040_168 0 0.008f
c211 id_M1_1040_248 0 0.008f
r106 id_M1_1040_248 id_M1_1040_252 0.4
c212 id_M1_1040_248 0 0.0004f
c213 id_M1_1040_252 0 0.0004f
r107 id_M1_1040_252 id_M1_1040_332 8.0
c214 id_M1_1040_252 0 0.008f
c215 id_M1_1040_332 0 0.008f
r108 id_M1_1040_332 id_M1_1040_412 8.0
c216 id_M1_1040_332 0 0.008f
c217 id_M1_1040_412 0 0.008f
r109 id_M1_1040_412 id_M1_1040_492 8.0
c218 id_M1_1040_412 0 0.008f
c219 id_M1_1040_492 0 0.008f
r110 id_M1_1040_492 id_M1_1040_504 1.2
c220 id_M1_1040_492 0 0.0012000000000000001f
c221 id_M1_1040_504 0 0.0012000000000000001f
r111 id_M1_1040_504 id_M1_1040_584 8.0
c222 id_M1_1040_504 0 0.008f
c223 id_M1_1040_584 0 0.008f
r112 id_M1_1040_584 id_M1_1040_664 8.0
c224 id_M1_1040_584 0 0.008f
c225 id_M1_1040_664 0 0.008f
r113 id_M1_1040_664 id_M1_1040_744 8.0
c226 id_M1_1040_664 0 0.008f
c227 id_M1_1040_744 0 0.008f
r114 id_M1_1040_744 id_M1_1040_792 4.8
c228 id_M1_1040_744 0 0.0048000000000000004f
c229 id_M1_1040_792 0 0.0048000000000000004f
r115 vss_M1_960_132 vss_M1_960_168 3.5999999999999996
c230 vss_M1_960_132 0 0.0036f
c231 vss_M1_960_168 0 0.0036f
r116 vss_M1_960_168 vss_M1_960_248 8.0
c232 vss_M1_960_168 0 0.008f
c233 vss_M1_960_248 0 0.008f
r117 vss_M1_960_248 vss_M1_960_328 8.0
c234 vss_M1_960_248 0 0.008f
c235 vss_M1_960_328 0 0.008f
r118 vss_M1_960_328 vss_M1_960_336 0.8
c236 vss_M1_960_328 0 0.0008f
c237 vss_M1_960_336 0 0.0008f
r119 vss_M1_960_336 vss_M1_960_416 8.0
c238 vss_M1_960_336 0 0.008f
c239 vss_M1_960_416 0 0.008f
r120 vss_M1_960_416 vss_M1_960_420 0.4
c240 vss_M1_960_416 0 0.0004f
c241 vss_M1_960_420 0 0.0004f
r121 vss_M1_960_420 vss_M1_960_462 4.2
c242 vss_M1_960_420 0 0.004200000000000001f
c243 vss_M1_960_462 0 0.004200000000000001f
r122 vss_M1_960_462 vss_M1_960_542 8.0
c244 vss_M1_960_462 0 0.008f
c245 vss_M1_960_542 0 0.008f
r123 vss_M1_960_542 vss_M1_960_588 4.6
c246 vss_M1_960_542 0 0.0046f
c247 vss_M1_960_588 0 0.0046f
r124 vss_M1_960_588 vss_M1_960_668 8.0
c248 vss_M1_960_588 0 0.008f
c249 vss_M1_960_668 0 0.008f
r125 vss_M1_960_668 vss_M1_960_748 8.0
c250 vss_M1_960_668 0 0.008f
c251 vss_M1_960_748 0 0.008f
r126 vss_M1_960_748 vss_M1_960_792 4.3999999999999995
c252 vss_M1_960_748 0 0.0044f
c253 vss_M1_960_792 0 0.0044f
r127 net10_M1_1120_132 net10_M1_1120_212 8.0
c254 net10_M1_1120_132 0 0.008f
c255 net10_M1_1120_212 0 0.008f
r128 net10_M1_1120_212 net10_M1_1120_292 8.0
c256 net10_M1_1120_212 0 0.008f
c257 net10_M1_1120_292 0 0.008f
r129 net10_M1_1120_292 net10_M1_1120_336 4.3999999999999995
c258 net10_M1_1120_292 0 0.0044f
c259 net10_M1_1120_336 0 0.0044f
r130 net10_M1_1120_336 net10_M1_1120_416 8.0
c260 net10_M1_1120_336 0 0.008f
c261 net10_M1_1120_416 0 0.008f
r131 net10_M1_1120_416 net10_M1_1120_462 4.6
c262 net10_M1_1120_416 0 0.0046f
c263 net10_M1_1120_462 0 0.0046f
r132 net10_M1_1120_462 net10_M1_1120_542 8.0
c264 net10_M1_1120_462 0 0.008f
c265 net10_M1_1120_542 0 0.008f
r133 net10_M1_1120_542 net10_M1_1120_588 4.6
c266 net10_M1_1120_542 0 0.0046f
c267 net10_M1_1120_588 0 0.0046f
r134 net10_M1_1120_588 net10_M1_1120_668 8.0
c268 net10_M1_1120_588 0 0.008f
c269 net10_M1_1120_668 0 0.008f
r135 net10_M1_1120_668 net10_M1_1120_748 8.0
c270 net10_M1_1120_668 0 0.008f
c271 net10_M1_1120_748 0 0.008f
r136 net10_M1_1120_748 net10_M1_1120_792 4.3999999999999995
c272 net10_M1_1120_748 0 0.0044f
c273 net10_M1_1120_792 0 0.0044f
r137 vinp_M1_1760_132 vinp_M1_1760_168 3.5999999999999996
c274 vinp_M1_1760_132 0 0.0036f
c275 vinp_M1_1760_168 0 0.0036f
r138 vinp_M1_1760_168 vinp_M1_1760_248 8.0
c276 vinp_M1_1760_168 0 0.008f
c277 vinp_M1_1760_248 0 0.008f
r139 vinp_M1_1760_248 vinp_M1_1760_328 8.0
c278 vinp_M1_1760_248 0 0.008f
c279 vinp_M1_1760_328 0 0.008f
r140 vinp_M1_1760_328 vinp_M1_1760_408 8.0
c280 vinp_M1_1760_328 0 0.008f
c281 vinp_M1_1760_408 0 0.008f
r141 vinp_M1_1760_408 vinp_M1_1760_420 1.2
c282 vinp_M1_1760_408 0 0.0012000000000000001f
c283 vinp_M1_1760_420 0 0.0012000000000000001f
r142 vinp_M1_1760_420 vinp_M1_1760_500 8.0
c284 vinp_M1_1760_420 0 0.008f
c285 vinp_M1_1760_500 0 0.008f
r143 vinp_M1_1760_500 vinp_M1_1760_580 8.0
c286 vinp_M1_1760_500 0 0.008f
c287 vinp_M1_1760_580 0 0.008f
r144 vinp_M1_1760_580 vinp_M1_1760_660 8.0
c288 vinp_M1_1760_580 0 0.008f
c289 vinp_M1_1760_660 0 0.008f
r145 vinp_M1_1760_660 vinp_M1_1760_740 8.0
c290 vinp_M1_1760_660 0 0.008f
c291 vinp_M1_1760_740 0 0.008f
r146 vinp_M1_1760_740 vinp_M1_1760_792 5.2
c292 vinp_M1_1760_740 0 0.0052f
c293 vinp_M1_1760_792 0 0.0052f
r147 net10_M1_1680_132 net10_M1_1680_168 3.5999999999999996
c294 net10_M1_1680_132 0 0.0036f
c295 net10_M1_1680_168 0 0.0036f
r148 net10_M1_1680_168 net10_M1_1680_248 8.0
c296 net10_M1_1680_168 0 0.008f
c297 net10_M1_1680_248 0 0.008f
r149 net10_M1_1680_248 net10_M1_1680_328 8.0
c298 net10_M1_1680_248 0 0.008f
c299 net10_M1_1680_328 0 0.008f
r150 net10_M1_1680_328 net10_M1_1680_336 0.8
c300 net10_M1_1680_328 0 0.0008f
c301 net10_M1_1680_336 0 0.0008f
r151 net10_M1_1680_336 net10_M1_1680_416 8.0
c302 net10_M1_1680_336 0 0.008f
c303 net10_M1_1680_416 0 0.008f
r152 net10_M1_1680_416 net10_M1_1680_462 4.6
c304 net10_M1_1680_416 0 0.0046f
c305 net10_M1_1680_462 0 0.0046f
r153 net10_M1_1680_462 net10_M1_1680_542 8.0
c306 net10_M1_1680_462 0 0.008f
c307 net10_M1_1680_542 0 0.008f
r154 net10_M1_1680_542 net10_M1_1680_588 4.6
c308 net10_M1_1680_542 0 0.0046f
c309 net10_M1_1680_588 0 0.0046f
r155 net10_M1_1680_588 net10_M1_1680_668 8.0
c310 net10_M1_1680_588 0 0.008f
c311 net10_M1_1680_668 0 0.008f
r156 net10_M1_1680_668 net10_M1_1680_748 8.0
c312 net10_M1_1680_668 0 0.008f
c313 net10_M1_1680_748 0 0.008f
r157 net10_M1_1680_748 net10_M1_1680_792 4.3999999999999995
c314 net10_M1_1680_748 0 0.0044f
c315 net10_M1_1680_792 0 0.0044f
r158 net8_M1_1840_132 net8_M1_1840_212 8.0
c316 net8_M1_1840_132 0 0.008f
c317 net8_M1_1840_212 0 0.008f
r159 net8_M1_1840_212 net8_M1_1840_252 4.0
c318 net8_M1_1840_212 0 0.004f
c319 net8_M1_1840_252 0 0.004f
r160 net8_M1_1840_252 net8_M1_1840_332 8.0
c320 net8_M1_1840_252 0 0.008f
c321 net8_M1_1840_332 0 0.008f
r161 net8_M1_1840_332 net8_M1_1840_336 0.4
c322 net8_M1_1840_332 0 0.0004f
c323 net8_M1_1840_336 0 0.0004f
r162 net8_M1_1840_336 net8_M1_1840_416 8.0
c324 net8_M1_1840_336 0 0.008f
c325 net8_M1_1840_416 0 0.008f
r163 net8_M1_1840_416 net8_M1_1840_462 4.6
c326 net8_M1_1840_416 0 0.0046f
c327 net8_M1_1840_462 0 0.0046f
r164 net8_M1_1840_462 net8_M1_1840_542 8.0
c328 net8_M1_1840_462 0 0.008f
c329 net8_M1_1840_542 0 0.008f
r165 net8_M1_1840_542 net8_M1_1840_588 4.6
c330 net8_M1_1840_542 0 0.0046f
c331 net8_M1_1840_588 0 0.0046f
r166 net8_M1_1840_588 net8_M1_1840_668 8.0
c332 net8_M1_1840_588 0 0.008f
c333 net8_M1_1840_668 0 0.008f
r167 net8_M1_1840_668 net8_M1_1840_748 8.0
c334 net8_M1_1840_668 0 0.008f
c335 net8_M1_1840_748 0 0.008f
r168 net8_M1_1840_748 net8_M1_1840_792 4.3999999999999995
c336 net8_M1_1840_748 0 0.0044f
c337 net8_M1_1840_792 0 0.0044f
r169 vinn_M1_2400_132 vinn_M1_2400_168 3.5999999999999996
c338 vinn_M1_2400_132 0 0.0036f
c339 vinn_M1_2400_168 0 0.0036f
r170 vinn_M1_2400_168 vinn_M1_2400_248 8.0
c340 vinn_M1_2400_168 0 0.008f
c341 vinn_M1_2400_248 0 0.008f
r171 vinn_M1_2400_248 vinn_M1_2400_328 8.0
c342 vinn_M1_2400_248 0 0.008f
c343 vinn_M1_2400_328 0 0.008f
r172 vinn_M1_2400_328 vinn_M1_2400_408 8.0
c344 vinn_M1_2400_328 0 0.008f
c345 vinn_M1_2400_408 0 0.008f
r173 vinn_M1_2400_408 vinn_M1_2400_488 8.0
c346 vinn_M1_2400_408 0 0.008f
c347 vinn_M1_2400_488 0 0.008f
r174 vinn_M1_2400_488 vinn_M1_2400_504 1.6
c348 vinn_M1_2400_488 0 0.0016f
c349 vinn_M1_2400_504 0 0.0016f
r175 vinn_M1_2400_504 vinn_M1_2400_584 8.0
c350 vinn_M1_2400_504 0 0.008f
c351 vinn_M1_2400_584 0 0.008f
r176 vinn_M1_2400_584 vinn_M1_2400_664 8.0
c352 vinn_M1_2400_584 0 0.008f
c353 vinn_M1_2400_664 0 0.008f
r177 vinn_M1_2400_664 vinn_M1_2400_744 8.0
c354 vinn_M1_2400_664 0 0.008f
c355 vinn_M1_2400_744 0 0.008f
r178 vinn_M1_2400_744 vinn_M1_2400_792 4.8
c356 vinn_M1_2400_744 0 0.0048000000000000004f
c357 vinn_M1_2400_792 0 0.0048000000000000004f
r179 net10_M1_2320_132 net10_M1_2320_168 3.5999999999999996
c358 net10_M1_2320_132 0 0.0036f
c359 net10_M1_2320_168 0 0.0036f
r180 net10_M1_2320_168 net10_M1_2320_248 8.0
c360 net10_M1_2320_168 0 0.008f
c361 net10_M1_2320_248 0 0.008f
r181 net10_M1_2320_248 net10_M1_2320_328 8.0
c362 net10_M1_2320_248 0 0.008f
c363 net10_M1_2320_328 0 0.008f
r182 net10_M1_2320_328 net10_M1_2320_336 0.8
c364 net10_M1_2320_328 0 0.0008f
c365 net10_M1_2320_336 0 0.0008f
r183 net10_M1_2320_336 net10_M1_2320_416 8.0
c366 net10_M1_2320_336 0 0.008f
c367 net10_M1_2320_416 0 0.008f
r184 net10_M1_2320_416 net10_M1_2320_462 4.6
c368 net10_M1_2320_416 0 0.0046f
c369 net10_M1_2320_462 0 0.0046f
r185 net10_M1_2320_462 net10_M1_2320_542 8.0
c370 net10_M1_2320_462 0 0.008f
c371 net10_M1_2320_542 0 0.008f
r186 net10_M1_2320_542 net10_M1_2320_588 4.6
c372 net10_M1_2320_542 0 0.0046f
c373 net10_M1_2320_588 0 0.0046f
r187 net10_M1_2320_588 net10_M1_2320_668 8.0
c374 net10_M1_2320_588 0 0.008f
c375 net10_M1_2320_668 0 0.008f
r188 net10_M1_2320_668 net10_M1_2320_748 8.0
c376 net10_M1_2320_668 0 0.008f
c377 net10_M1_2320_748 0 0.008f
r189 net10_M1_2320_748 net10_M1_2320_792 4.3999999999999995
c378 net10_M1_2320_748 0 0.0044f
c379 net10_M1_2320_792 0 0.0044f
r190 vout_M1_2480_132 vout_M1_2480_212 8.0
c380 vout_M1_2480_132 0 0.008f
c381 vout_M1_2480_212 0 0.008f
r191 vout_M1_2480_212 vout_M1_2480_292 8.0
c382 vout_M1_2480_212 0 0.008f
c383 vout_M1_2480_292 0 0.008f
r192 vout_M1_2480_292 vout_M1_2480_336 4.3999999999999995
c384 vout_M1_2480_292 0 0.0044f
c385 vout_M1_2480_336 0 0.0044f
r193 vout_M1_2480_336 vout_M1_2480_416 8.0
c386 vout_M1_2480_336 0 0.008f
c387 vout_M1_2480_416 0 0.008f
r194 vout_M1_2480_416 vout_M1_2480_462 4.6
c388 vout_M1_2480_416 0 0.0046f
c389 vout_M1_2480_462 0 0.0046f
r195 vout_M1_2480_462 vout_M1_2480_542 8.0
c390 vout_M1_2480_462 0 0.008f
c391 vout_M1_2480_542 0 0.008f
r196 vout_M1_2480_542 vout_M1_2480_588 4.6
c392 vout_M1_2480_542 0 0.0046f
c393 vout_M1_2480_588 0 0.0046f
r197 vout_M1_2480_588 vout_M1_2480_668 8.0
c394 vout_M1_2480_588 0 0.008f
c395 vout_M1_2480_668 0 0.008f
r198 vout_M1_2480_668 vout_M1_2480_748 8.0
c396 vout_M1_2480_668 0 0.008f
c397 vout_M1_2480_748 0 0.008f
r199 vout_M1_2480_748 vout_M1_2480_792 4.3999999999999995
c398 vout_M1_2480_748 0 0.0044f
c399 vout_M1_2480_792 0 0.0044f
r200 vss_M2_284_168 vss_M2_320_168 2.1599999999999997
c400 vss_M2_284_168 0 0.0036f
c401 vss_M2_320_168 0 0.0036f
r201 vss_M2_320_168 vss_M2_400_168 4.8
c402 vss_M2_320_168 0 0.008f
c403 vss_M2_400_168 0 0.008f
r202 vss_M2_400_168 vss_M2_480_168 4.8
c404 vss_M2_400_168 0 0.008f
c405 vss_M2_480_168 0 0.008f
r203 vss_M2_480_168 vss_M2_560_168 4.8
c406 vss_M2_480_168 0 0.008f
c407 vss_M2_560_168 0 0.008f
r204 vss_M2_560_168 vss_M2_640_168 4.8
c408 vss_M2_560_168 0 0.008f
c409 vss_M2_640_168 0 0.008f
r205 vss_M2_640_168 vss_M2_720_168 4.8
c410 vss_M2_640_168 0 0.008f
c411 vss_M2_720_168 0 0.008f
r206 vss_M2_720_168 vss_M2_800_168 4.8
c412 vss_M2_720_168 0 0.008f
c413 vss_M2_800_168 0 0.008f
r207 vss_M2_800_168 vss_M2_880_168 4.8
c414 vss_M2_800_168 0 0.008f
c415 vss_M2_880_168 0 0.008f
r208 vss_M2_880_168 vss_M2_960_168 4.8
c416 vss_M2_880_168 0 0.008f
c417 vss_M2_960_168 0 0.008f
r209 vss_M2_960_168 vss_M2_996_168 2.1599999999999997
c418 vss_M2_960_168 0 0.0036f
c419 vss_M2_996_168 0 0.0036f
r210 net10_M2_1244_168 net10_M2_1280_168 2.1599999999999997
c420 net10_M2_1244_168 0 0.0036f
c421 net10_M2_1280_168 0 0.0036f
r211 net10_M2_1280_168 net10_M2_1360_168 4.8
c422 net10_M2_1280_168 0 0.008f
c423 net10_M2_1360_168 0 0.008f
r212 net10_M2_1360_168 net10_M2_1440_168 4.8
c424 net10_M2_1360_168 0 0.008f
c425 net10_M2_1440_168 0 0.008f
r213 net10_M2_1440_168 net10_M2_1520_168 4.8
c426 net10_M2_1440_168 0 0.008f
c427 net10_M2_1520_168 0 0.008f
r214 net10_M2_1520_168 net10_M2_1600_168 4.8
c428 net10_M2_1520_168 0 0.008f
c429 net10_M2_1600_168 0 0.008f
r215 net10_M2_1600_168 net10_M2_1680_168 4.8
c430 net10_M2_1600_168 0 0.008f
c431 net10_M2_1680_168 0 0.008f
r216 net10_M2_1680_168 net10_M2_1760_168 4.8
c432 net10_M2_1680_168 0 0.008f
c433 net10_M2_1760_168 0 0.008f
r217 net10_M2_1760_168 net10_M2_1840_168 4.8
c434 net10_M2_1760_168 0 0.008f
c435 net10_M2_1840_168 0 0.008f
r218 net10_M2_1840_168 net10_M2_1920_168 4.8
c436 net10_M2_1840_168 0 0.008f
c437 net10_M2_1920_168 0 0.008f
r219 net10_M2_1920_168 net10_M2_2000_168 4.8
c438 net10_M2_1920_168 0 0.008f
c439 net10_M2_2000_168 0 0.008f
r220 net10_M2_2000_168 net10_M2_2080_168 4.8
c440 net10_M2_2000_168 0 0.008f
c441 net10_M2_2080_168 0 0.008f
r221 net10_M2_2080_168 net10_M2_2160_168 4.8
c442 net10_M2_2080_168 0 0.008f
c443 net10_M2_2160_168 0 0.008f
r222 net10_M2_2160_168 net10_M2_2240_168 4.8
c444 net10_M2_2160_168 0 0.008f
c445 net10_M2_2240_168 0 0.008f
r223 net10_M2_2240_168 net10_M2_2320_168 4.8
c446 net10_M2_2240_168 0 0.008f
c447 net10_M2_2320_168 0 0.008f
r224 net10_M2_2320_168 net10_M2_2356_168 2.1599999999999997
c448 net10_M2_2320_168 0 0.0036f
c449 net10_M2_2356_168 0 0.0036f
r225 vdd_M2_3004_168 vdd_M2_3040_168 2.1599999999999997
c450 vdd_M2_3004_168 0 0.0036f
c451 vdd_M2_3040_168 0 0.0036f
r226 vdd_M2_3040_168 vdd_M2_3120_168 4.8
c452 vdd_M2_3040_168 0 0.008f
c453 vdd_M2_3120_168 0 0.008f
r227 vdd_M2_3120_168 vdd_M2_3200_168 4.8
c454 vdd_M2_3120_168 0 0.008f
c455 vdd_M2_3200_168 0 0.008f
r228 vdd_M2_3200_168 vdd_M2_3280_168 4.8
c456 vdd_M2_3200_168 0 0.008f
c457 vdd_M2_3280_168 0 0.008f
r229 vdd_M2_3280_168 vdd_M2_3316_168 2.1599999999999997
c458 vdd_M2_3280_168 0 0.0036f
c459 vdd_M2_3316_168 0 0.0036f
r230 vdd_M2_3724_168 vdd_M2_3760_168 2.1599999999999997
c460 vdd_M2_3724_168 0 0.0036f
c461 vdd_M2_3760_168 0 0.0036f
r231 vdd_M2_3760_168 vdd_M2_3840_168 4.8
c462 vdd_M2_3760_168 0 0.008f
c463 vdd_M2_3840_168 0 0.008f
r232 vdd_M2_3840_168 vdd_M2_3920_168 4.8
c464 vdd_M2_3840_168 0 0.008f
c465 vdd_M2_3920_168 0 0.008f
r233 vdd_M2_3920_168 vdd_M2_3956_168 2.1599999999999997
c466 vdd_M2_3920_168 0 0.0036f
c467 vdd_M2_3956_168 0 0.0036f
r234 net10_M2_684_336 net10_M2_720_336 2.1599999999999997
c468 net10_M2_684_336 0 0.0036f
c469 net10_M2_720_336 0 0.0036f
r235 net10_M2_720_336 net10_M2_800_336 4.8
c470 net10_M2_720_336 0 0.008f
c471 net10_M2_800_336 0 0.008f
r236 net10_M2_800_336 net10_M2_880_336 4.8
c472 net10_M2_800_336 0 0.008f
c473 net10_M2_880_336 0 0.008f
r237 net10_M2_880_336 net10_M2_960_336 4.8
c474 net10_M2_880_336 0 0.008f
c475 net10_M2_960_336 0 0.008f
r238 net10_M2_960_336 net10_M2_1040_336 4.8
c476 net10_M2_960_336 0 0.008f
c477 net10_M2_1040_336 0 0.008f
r239 net10_M2_1040_336 net10_M2_1120_336 4.8
c478 net10_M2_1040_336 0 0.008f
c479 net10_M2_1120_336 0 0.008f
r240 net10_M2_1120_336 net10_M2_1156_336 2.1599999999999997
c480 net10_M2_1120_336 0 0.0036f
c481 net10_M2_1156_336 0 0.0036f
r241 vout_M2_2284_336 vout_M2_2364_336 4.8
c482 vout_M2_2284_336 0 0.008f
c483 vout_M2_2364_336 0 0.008f
r242 vout_M2_2364_336 vout_M2_2444_336 4.8
c484 vout_M2_2364_336 0 0.008f
c485 vout_M2_2444_336 0 0.008f
r243 vout_M2_2444_336 vout_M2_2480_336 2.1599999999999997
c486 vout_M2_2444_336 0 0.0036f
c487 vout_M2_2480_336 0 0.0036f
r244 vout_M2_2480_336 vout_M2_2560_336 4.8
c488 vout_M2_2480_336 0 0.008f
c489 vout_M2_2560_336 0 0.008f
r245 vout_M2_2560_336 vout_M2_2580_336 1.2
c490 vout_M2_2560_336 0 0.002f
c491 vout_M2_2580_336 0 0.002f
r246 net8_M2_2844_336 net8_M2_2880_336 2.1599999999999997
c492 net8_M2_2844_336 0 0.0036f
c493 net8_M2_2880_336 0 0.0036f
r247 net8_M2_2880_336 net8_M2_2960_336 4.8
c494 net8_M2_2880_336 0 0.008f
c495 net8_M2_2960_336 0 0.008f
r248 net8_M2_2960_336 net8_M2_3040_336 4.8
c496 net8_M2_2960_336 0 0.008f
c497 net8_M2_3040_336 0 0.008f
r249 net8_M2_3040_336 net8_M2_3120_336 4.8
c498 net8_M2_3040_336 0 0.008f
c499 net8_M2_3120_336 0 0.008f
r250 net8_M2_3120_336 net8_M2_3200_336 4.8
c500 net8_M2_3120_336 0 0.008f
c501 net8_M2_3200_336 0 0.008f
r251 net8_M2_3200_336 net8_M2_3236_336 2.1599999999999997
c502 net8_M2_3200_336 0 0.0036f
c503 net8_M2_3236_336 0 0.0036f
r252 vdd_M2_3324_336 vdd_M2_3360_336 2.1599999999999997
c504 vdd_M2_3324_336 0 0.0036f
c505 vdd_M2_3360_336 0 0.0036f
r253 vdd_M2_3360_336 vdd_M2_3440_336 4.8
c506 vdd_M2_3360_336 0 0.008f
c507 vdd_M2_3440_336 0 0.008f
r254 vdd_M2_3440_336 vdd_M2_3520_336 4.8
c508 vdd_M2_3440_336 0 0.008f
c509 vdd_M2_3520_336 0 0.008f
r255 vdd_M2_3520_336 vdd_M2_3600_336 4.8
c510 vdd_M2_3520_336 0 0.008f
c511 vdd_M2_3600_336 0 0.008f
r256 vdd_M2_3600_336 vdd_M2_3636_336 2.1599999999999997
c512 vdd_M2_3600_336 0 0.0036f
c513 vdd_M2_3636_336 0 0.0036f
r257 vdd_M2_3724_336 vdd_M2_3760_336 2.1599999999999997
c514 vdd_M2_3724_336 0 0.0036f
c515 vdd_M2_3760_336 0 0.0036f
r258 vdd_M2_3760_336 vdd_M2_3840_336 4.8
c516 vdd_M2_3760_336 0 0.008f
c517 vdd_M2_3840_336 0 0.008f
r259 vdd_M2_3840_336 vdd_M2_3920_336 4.8
c518 vdd_M2_3840_336 0 0.008f
c519 vdd_M2_3920_336 0 0.008f
r260 vdd_M2_3920_336 vdd_M2_3956_336 2.1599999999999997
c520 vdd_M2_3920_336 0 0.0036f
c521 vdd_M2_3956_336 0 0.0036f
r261 id_M2_364_252 id_M2_400_252 2.1599999999999997
c522 id_M2_364_252 0 0.0036f
c523 id_M2_400_252 0 0.0036f
r262 id_M2_400_252 id_M2_480_252 4.8
c524 id_M2_400_252 0 0.008f
c525 id_M2_480_252 0 0.008f
r263 id_M2_480_252 id_M2_560_252 4.8
c526 id_M2_480_252 0 0.008f
c527 id_M2_560_252 0 0.008f
r264 id_M2_560_252 id_M2_640_252 4.8
c528 id_M2_560_252 0 0.008f
c529 id_M2_640_252 0 0.008f
r265 id_M2_640_252 id_M2_720_252 4.8
c530 id_M2_640_252 0 0.008f
c531 id_M2_720_252 0 0.008f
r266 id_M2_720_252 id_M2_800_252 4.8
c532 id_M2_720_252 0 0.008f
c533 id_M2_800_252 0 0.008f
r267 id_M2_800_252 id_M2_880_252 4.8
c534 id_M2_800_252 0 0.008f
c535 id_M2_880_252 0 0.008f
r268 id_M2_880_252 id_M2_960_252 4.8
c536 id_M2_880_252 0 0.008f
c537 id_M2_960_252 0 0.008f
r269 id_M2_960_252 id_M2_1040_252 4.8
c538 id_M2_960_252 0 0.008f
c539 id_M2_1040_252 0 0.008f
r270 id_M2_1040_252 id_M2_1076_252 2.1599999999999997
c540 id_M2_1040_252 0 0.0036f
c541 id_M2_1076_252 0 0.0036f
r271 vinp_M2_1324_252 vinp_M2_1360_252 2.1599999999999997
c542 vinp_M2_1324_252 0 0.0036f
c543 vinp_M2_1360_252 0 0.0036f
r272 vinp_M2_1360_252 vinp_M2_1440_252 4.8
c544 vinp_M2_1360_252 0 0.008f
c545 vinp_M2_1440_252 0 0.008f
r273 vinp_M2_1440_252 vinp_M2_1520_252 4.8
c546 vinp_M2_1440_252 0 0.008f
c547 vinp_M2_1520_252 0 0.008f
r274 vinp_M2_1520_252 vinp_M2_1600_252 4.8
c548 vinp_M2_1520_252 0 0.008f
c549 vinp_M2_1600_252 0 0.008f
r275 vinp_M2_1600_252 vinp_M2_1636_252 2.1599999999999997
c550 vinp_M2_1600_252 0 0.0036f
c551 vinp_M2_1636_252 0 0.0036f
r276 net8_M2_1804_252 net8_M2_1840_252 2.1599999999999997
c552 net8_M2_1804_252 0 0.0036f
c553 net8_M2_1840_252 0 0.0036f
r277 net8_M2_1840_252 net8_M2_1920_252 4.8
c554 net8_M2_1840_252 0 0.008f
c555 net8_M2_1920_252 0 0.008f
r278 net8_M2_1920_252 net8_M2_2000_252 4.8
c556 net8_M2_1920_252 0 0.008f
c557 net8_M2_2000_252 0 0.008f
r279 net8_M2_2000_252 net8_M2_2080_252 4.8
c558 net8_M2_2000_252 0 0.008f
c559 net8_M2_2080_252 0 0.008f
r280 net8_M2_2080_252 net8_M2_2160_252 4.8
c560 net8_M2_2080_252 0 0.008f
c561 net8_M2_2160_252 0 0.008f
r281 net8_M2_2160_252 net8_M2_2196_252 2.1599999999999997
c562 net8_M2_2160_252 0 0.0036f
c563 net8_M2_2196_252 0 0.0036f
r282 vout_M2_2364_252 vout_M2_2400_252 2.1599999999999997
c564 vout_M2_2364_252 0 0.0036f
c565 vout_M2_2400_252 0 0.0036f
r283 vout_M2_2400_252 vout_M2_2480_252 4.8
c566 vout_M2_2400_252 0 0.008f
c567 vout_M2_2480_252 0 0.008f
r284 vout_M2_2480_252 vout_M2_2560_252 4.8
c568 vout_M2_2480_252 0 0.008f
c569 vout_M2_2560_252 0 0.008f
r285 vout_M2_2560_252 vout_M2_2640_252 4.8
c570 vout_M2_2560_252 0 0.008f
c571 vout_M2_2640_252 0 0.008f
r286 vout_M2_2640_252 vout_M2_2676_252 2.1599999999999997
c572 vout_M2_2640_252 0 0.0036f
c573 vout_M2_2676_252 0 0.0036f
r287 vout_M2_2924_252 vout_M2_2960_252 2.1599999999999997
c574 vout_M2_2924_252 0 0.0036f
c575 vout_M2_2960_252 0 0.0036f
r288 vout_M2_2960_252 vout_M2_3040_252 4.8
c576 vout_M2_2960_252 0 0.008f
c577 vout_M2_3040_252 0 0.008f
r289 vout_M2_3040_252 vout_M2_3120_252 4.8
c578 vout_M2_3040_252 0 0.008f
c579 vout_M2_3120_252 0 0.008f
r290 vout_M2_3120_252 vout_M2_3200_252 4.8
c580 vout_M2_3120_252 0 0.008f
c581 vout_M2_3200_252 0 0.008f
r291 vout_M2_3200_252 vout_M2_3236_252 2.1599999999999997
c582 vout_M2_3200_252 0 0.0036f
c583 vout_M2_3236_252 0 0.0036f
r292 net8_M2_3644_252 net8_M2_3680_252 2.1599999999999997
c584 net8_M2_3644_252 0 0.0036f
c585 net8_M2_3680_252 0 0.0036f
r293 net8_M2_3680_252 net8_M2_3760_252 4.8
c586 net8_M2_3680_252 0 0.008f
c587 net8_M2_3760_252 0 0.008f
r294 net8_M2_3760_252 net8_M2_3840_252 4.8
c588 net8_M2_3760_252 0 0.008f
c589 net8_M2_3840_252 0 0.008f
r295 net8_M2_3840_252 net8_M2_3920_252 4.8
c590 net8_M2_3840_252 0 0.008f
c591 net8_M2_3920_252 0 0.008f
r296 net8_M2_3920_252 net8_M2_3956_252 2.1599999999999997
c592 net8_M2_3920_252 0 0.0036f
c593 net8_M2_3956_252 0 0.0036f
r297 vss_M2_284_420 vss_M2_320_420 2.1599999999999997
c594 vss_M2_284_420 0 0.0036f
c595 vss_M2_320_420 0 0.0036f
r298 vss_M2_320_420 vss_M2_400_420 4.8
c596 vss_M2_320_420 0 0.008f
c597 vss_M2_400_420 0 0.008f
r299 vss_M2_400_420 vss_M2_480_420 4.8
c598 vss_M2_400_420 0 0.008f
c599 vss_M2_480_420 0 0.008f
r300 vss_M2_480_420 vss_M2_560_420 4.8
c600 vss_M2_480_420 0 0.008f
c601 vss_M2_560_420 0 0.008f
r301 vss_M2_560_420 vss_M2_640_420 4.8
c602 vss_M2_560_420 0 0.008f
c603 vss_M2_640_420 0 0.008f
r302 vss_M2_640_420 vss_M2_720_420 4.8
c604 vss_M2_640_420 0 0.008f
c605 vss_M2_720_420 0 0.008f
r303 vss_M2_720_420 vss_M2_800_420 4.8
c606 vss_M2_720_420 0 0.008f
c607 vss_M2_800_420 0 0.008f
r304 vss_M2_800_420 vss_M2_880_420 4.8
c608 vss_M2_800_420 0 0.008f
c609 vss_M2_880_420 0 0.008f
r305 vss_M2_880_420 vss_M2_960_420 4.8
c610 vss_M2_880_420 0 0.008f
c611 vss_M2_960_420 0 0.008f
r306 vss_M2_960_420 vss_M2_996_420 2.1599999999999997
c612 vss_M2_960_420 0 0.0036f
c613 vss_M2_996_420 0 0.0036f
r307 vinp_M2_1724_420 vinp_M2_1760_420 2.1599999999999997
c614 vinp_M2_1724_420 0 0.0036f
c615 vinp_M2_1760_420 0 0.0036f
r308 vinp_M2_1760_420 vinp_M2_1840_420 4.8
c616 vinp_M2_1760_420 0 0.008f
c617 vinp_M2_1840_420 0 0.008f
r309 vinp_M2_1840_420 vinp_M2_1920_420 4.8
c618 vinp_M2_1840_420 0 0.008f
c619 vinp_M2_1920_420 0 0.008f
r310 vinp_M2_1920_420 vinp_M2_2000_420 4.8
c620 vinp_M2_1920_420 0 0.008f
c621 vinp_M2_2000_420 0 0.008f
r311 vinp_M2_2000_420 vinp_M2_2020_420 1.2
c622 vinp_M2_2000_420 0 0.002f
c623 vinp_M2_2020_420 0 0.002f
r312 vdd_M2_3004_420 vdd_M2_3040_420 2.1599999999999997
c624 vdd_M2_3004_420 0 0.0036f
c625 vdd_M2_3040_420 0 0.0036f
r313 vdd_M2_3040_420 vdd_M2_3120_420 4.8
c626 vdd_M2_3040_420 0 0.008f
c627 vdd_M2_3120_420 0 0.008f
r314 vdd_M2_3120_420 vdd_M2_3200_420 4.8
c628 vdd_M2_3120_420 0 0.008f
c629 vdd_M2_3200_420 0 0.008f
r315 vdd_M2_3200_420 vdd_M2_3280_420 4.8
c630 vdd_M2_3200_420 0 0.008f
c631 vdd_M2_3280_420 0 0.008f
r316 vdd_M2_3280_420 vdd_M2_3316_420 2.1599999999999997
c632 vdd_M2_3280_420 0 0.0036f
c633 vdd_M2_3316_420 0 0.0036f
r317 net8_M2_3644_420 net8_M2_3680_420 2.1599999999999997
c634 net8_M2_3644_420 0 0.0036f
c635 net8_M2_3680_420 0 0.0036f
r318 net8_M2_3680_420 net8_M2_3760_420 4.8
c636 net8_M2_3680_420 0 0.008f
c637 net8_M2_3760_420 0 0.008f
r319 net8_M2_3760_420 net8_M2_3840_420 4.8
c638 net8_M2_3760_420 0 0.008f
c639 net8_M2_3840_420 0 0.008f
r320 net8_M2_3840_420 net8_M2_3920_420 4.8
c640 net8_M2_3840_420 0 0.008f
c641 net8_M2_3920_420 0 0.008f
r321 net8_M2_3920_420 net8_M2_3956_420 2.1599999999999997
c642 net8_M2_3920_420 0 0.0036f
c643 net8_M2_3956_420 0 0.0036f
r322 id_M2_364_504 id_M2_400_504 2.1599999999999997
c644 id_M2_364_504 0 0.0036f
c645 id_M2_400_504 0 0.0036f
r323 id_M2_400_504 id_M2_480_504 4.8
c646 id_M2_400_504 0 0.008f
c647 id_M2_480_504 0 0.008f
r324 id_M2_480_504 id_M2_560_504 4.8
c648 id_M2_480_504 0 0.008f
c649 id_M2_560_504 0 0.008f
r325 id_M2_560_504 id_M2_640_504 4.8
c650 id_M2_560_504 0 0.008f
c651 id_M2_640_504 0 0.008f
r326 id_M2_640_504 id_M2_720_504 4.8
c652 id_M2_640_504 0 0.008f
c653 id_M2_720_504 0 0.008f
r327 id_M2_720_504 id_M2_800_504 4.8
c654 id_M2_720_504 0 0.008f
c655 id_M2_800_504 0 0.008f
r328 id_M2_800_504 id_M2_880_504 4.8
c656 id_M2_800_504 0 0.008f
c657 id_M2_880_504 0 0.008f
r329 id_M2_880_504 id_M2_960_504 4.8
c658 id_M2_880_504 0 0.008f
c659 id_M2_960_504 0 0.008f
r330 id_M2_960_504 id_M2_1040_504 4.8
c660 id_M2_960_504 0 0.008f
c661 id_M2_1040_504 0 0.008f
r331 id_M2_1040_504 id_M2_1076_504 2.1599999999999997
c662 id_M2_1040_504 0 0.0036f
c663 id_M2_1076_504 0 0.0036f
r332 vinn_M2_2204_504 vinn_M2_2284_504 4.8
c664 vinn_M2_2204_504 0 0.008f
c665 vinn_M2_2284_504 0 0.008f
r333 vinn_M2_2284_504 vinn_M2_2364_504 4.8
c666 vinn_M2_2284_504 0 0.008f
c667 vinn_M2_2364_504 0 0.008f
r334 vinn_M2_2364_504 vinn_M2_2400_504 2.1599999999999997
c668 vinn_M2_2364_504 0 0.0036f
c669 vinn_M2_2400_504 0 0.0036f
r335 vinn_M2_2400_504 vinn_M2_2436_504 2.1599999999999997
c670 vinn_M2_2400_504 0 0.0036f
c671 vinn_M2_2436_504 0 0.0036f
r336 vout_M2_2924_504 vout_M2_2960_504 2.1599999999999997
c672 vout_M2_2924_504 0 0.0036f
c673 vout_M2_2960_504 0 0.0036f
r337 vout_M2_2960_504 vout_M2_3040_504 4.8
c674 vout_M2_2960_504 0 0.008f
c675 vout_M2_3040_504 0 0.008f
r338 vout_M2_3040_504 vout_M2_3120_504 4.8
c676 vout_M2_3040_504 0 0.008f
c677 vout_M2_3120_504 0 0.008f
r339 vout_M2_3120_504 vout_M2_3200_504 4.8
c678 vout_M2_3120_504 0 0.008f
c679 vout_M2_3200_504 0 0.008f
r340 vout_M2_3200_504 vout_M2_3236_504 2.1599999999999997
c680 vout_M2_3200_504 0 0.0036f
c681 vout_M2_3236_504 0 0.0036f
r341 net10_M2_684_588 net10_M2_720_588 2.1599999999999997
c682 net10_M2_684_588 0 0.0036f
c683 net10_M2_720_588 0 0.0036f
r342 net10_M2_720_588 net10_M2_800_588 4.8
c684 net10_M2_720_588 0 0.008f
c685 net10_M2_800_588 0 0.008f
r343 net10_M2_800_588 net10_M2_880_588 4.8
c686 net10_M2_800_588 0 0.008f
c687 net10_M2_880_588 0 0.008f
r344 net10_M2_880_588 net10_M2_960_588 4.8
c688 net10_M2_880_588 0 0.008f
c689 net10_M2_960_588 0 0.008f
r345 net10_M2_960_588 net10_M2_1040_588 4.8
c690 net10_M2_960_588 0 0.008f
c691 net10_M2_1040_588 0 0.008f
r346 net10_M2_1040_588 net10_M2_1120_588 4.8
c692 net10_M2_1040_588 0 0.008f
c693 net10_M2_1120_588 0 0.008f
r347 net10_M2_1120_588 net10_M2_1156_588 2.1599999999999997
c694 net10_M2_1120_588 0 0.0036f
c695 net10_M2_1156_588 0 0.0036f
r348 net8_M2_2844_588 net8_M2_2880_588 2.1599999999999997
c696 net8_M2_2844_588 0 0.0036f
c697 net8_M2_2880_588 0 0.0036f
r349 net8_M2_2880_588 net8_M2_2960_588 4.8
c698 net8_M2_2880_588 0 0.008f
c699 net8_M2_2960_588 0 0.008f
r350 net8_M2_2960_588 net8_M2_3040_588 4.8
c700 net8_M2_2960_588 0 0.008f
c701 net8_M2_3040_588 0 0.008f
r351 net8_M2_3040_588 net8_M2_3120_588 4.8
c702 net8_M2_3040_588 0 0.008f
c703 net8_M2_3120_588 0 0.008f
r352 net8_M2_3120_588 net8_M2_3200_588 4.8
c704 net8_M2_3120_588 0 0.008f
c705 net8_M2_3200_588 0 0.008f
r353 net8_M2_3200_588 net8_M2_3236_588 2.1599999999999997
c706 net8_M2_3200_588 0 0.0036f
c707 net8_M2_3236_588 0 0.0036f
r354 id_M2_540_0 id_M2_620_0 4.8
c708 id_M2_540_0 0 0.008f
c709 id_M2_620_0 0 0.008f
r355 id_M2_620_0 id_M2_640_0 1.2
c710 id_M2_620_0 0 0.002f
c711 id_M2_640_0 0 0.002f
r356 id_M2_640_0 id_M2_720_0 4.8
c712 id_M2_640_0 0 0.008f
c713 id_M2_720_0 0 0.008f
r357 id_M2_720_0 id_M2_740_0 1.2
c714 id_M2_720_0 0 0.002f
c715 id_M2_740_0 0 0.002f
r358 vinp_M2_1324_0 vinp_M2_1360_0 2.1599999999999997
c716 vinp_M2_1324_0 0 0.0036f
c717 vinp_M2_1360_0 0 0.0036f
r359 vinp_M2_1360_0 vinp_M2_1440_0 4.8
c718 vinp_M2_1360_0 0 0.008f
c719 vinp_M2_1440_0 0 0.008f
r360 vinp_M2_1440_0 vinp_M2_1520_0 4.8
c720 vinp_M2_1440_0 0 0.008f
c721 vinp_M2_1520_0 0 0.008f
r361 vinp_M2_1520_0 vinp_M2_1600_0 4.8
c722 vinp_M2_1520_0 0 0.008f
c723 vinp_M2_1600_0 0 0.008f
r362 vinp_M2_1600_0 vinp_M2_1680_0 4.8
c724 vinp_M2_1600_0 0 0.008f
c725 vinp_M2_1680_0 0 0.008f
r363 vinp_M2_1680_0 vinp_M2_1760_0 4.8
c726 vinp_M2_1680_0 0 0.008f
c727 vinp_M2_1760_0 0 0.008f
r364 vinp_M2_1760_0 vinp_M2_1840_0 4.8
c728 vinp_M2_1760_0 0 0.008f
c729 vinp_M2_1840_0 0 0.008f
r365 vout_M2_2300_0 vout_M2_2380_0 4.8
c730 vout_M2_2300_0 0 0.008f
c731 vout_M2_2380_0 0 0.008f
r366 vout_M2_2380_0 vout_M2_2400_0 1.2
c732 vout_M2_2380_0 0 0.002f
c733 vout_M2_2400_0 0 0.002f
r367 vout_M2_2400_0 vout_M2_2480_0 4.8
c734 vout_M2_2400_0 0 0.008f
c735 vout_M2_2480_0 0 0.008f
r368 vout_M2_2480_0 vout_M2_2500_0 1.2
c736 vout_M2_2480_0 0 0.002f
c737 vout_M2_2500_0 0 0.002f
r369 vdd_M2_3820_0 vdd_M2_3900_0 4.8
c738 vdd_M2_3820_0 0 0.008f
c739 vdd_M2_3900_0 0 0.008f
r370 vdd_M2_3900_0 vdd_M2_3920_0 1.2
c740 vdd_M2_3900_0 0 0.002f
c741 vdd_M2_3920_0 0 0.002f
r371 vdd_M2_3920_0 vdd_M2_4000_0 4.8
c742 vdd_M2_3920_0 0 0.008f
c743 vdd_M2_4000_0 0 0.008f
r372 vdd_M2_4000_0 vdd_M2_4020_0 1.2
c744 vdd_M2_4000_0 0 0.002f
c745 vdd_M2_4020_0 0 0.002f
r373 vout_M2_2444_84 vout_M2_2480_84 2.1599999999999997
c746 vout_M2_2444_84 0 0.0036f
c747 vout_M2_2480_84 0 0.0036f
r374 vout_M2_2480_84 vout_M2_2560_84 4.8
c748 vout_M2_2480_84 0 0.008f
c749 vout_M2_2560_84 0 0.008f
r375 vout_M2_2560_84 vout_M2_2640_84 4.8
c750 vout_M2_2560_84 0 0.008f
c751 vout_M2_2640_84 0 0.008f
r376 vout_M2_2640_84 vout_M2_2720_84 4.8
c752 vout_M2_2640_84 0 0.008f
c753 vout_M2_2720_84 0 0.008f
r377 vout_M2_2720_84 vout_M2_2800_84 4.8
c754 vout_M2_2720_84 0 0.008f
c755 vout_M2_2800_84 0 0.008f
r378 vout_M2_2800_84 vout_M2_2880_84 4.8
c756 vout_M2_2800_84 0 0.008f
c757 vout_M2_2880_84 0 0.008f
r379 vout_M2_2880_84 vout_M2_2960_84 4.8
c758 vout_M2_2880_84 0 0.008f
c759 vout_M2_2960_84 0 0.008f
r380 vout_M2_2960_84 vout_M2_2996_84 2.1599999999999997
c760 vout_M2_2960_84 0 0.0036f
c761 vout_M2_2996_84 0 0.0036f
r381 vdd_M1_3920_168 vdd_M2_3920_168 50
r382 vdd_M1_3920_336 vdd_M2_3920_336 50
r383 net8_M1_3840_252 net8_M2_3840_252 50
r384 net8_M1_3840_420 net8_M2_3840_420 50
r385 net8_M1_3760_252 net8_M2_3760_252 50
r386 net8_M1_3760_420 net8_M2_3760_420 50
r387 vdd_M1_3200_168 vdd_M2_3200_168 50
r388 vdd_M1_3200_420 vdd_M2_3200_420 50
r389 vout_M1_3040_252 vout_M2_3040_252 50
r390 vout_M1_3040_504 vout_M2_3040_504 50
r391 net8_M1_3120_336 net8_M2_3120_336 50
r392 net8_M1_3120_588 net8_M2_3120_588 50
r393 vss_M1_960_168 vss_M2_960_168 50
r394 vss_M1_960_420 vss_M2_960_420 50
r395 vss_M1_320_168 vss_M2_320_168 50
r396 vss_M1_320_420 vss_M2_320_420 50
r397 id_M1_1040_252 id_M2_1040_252 50
r398 id_M1_1040_504 id_M2_1040_504 50
r399 id_M1_400_252 id_M2_400_252 50
r400 id_M1_400_504 id_M2_400_504 50
r401 id_M1_480_252 id_M2_480_252 50
r402 id_M1_480_504 id_M2_480_504 50
r403 net10_M1_1120_336 net10_M2_1120_336 50
r404 net10_M1_1120_588 net10_M2_1120_588 50
r405 net10_M1_2320_168 net10_M2_2320_168 50
r406 net10_M1_1680_168 net10_M2_1680_168 50
r407 net8_M1_1840_252 net8_M2_1840_252 50
r408 vout_M1_2480_336 vout_M2_2480_336 50
r409 vinp_M1_1760_420 vinp_M2_1760_420 50
r410 vinn_M1_2400_504 vinn_M2_2400_504 50
r411 vdd_M3_3920__36 vdd_M3_3920_0 1.44
c762 vdd_M3_3920__36 0 0.0036f
c763 vdd_M3_3920_0 0 0.0036f
r412 vdd_M3_3920_0 vdd_M3_3920_80 3.2
c764 vdd_M3_3920_0 0 0.008f
c765 vdd_M3_3920_80 0 0.008f
r413 vdd_M3_3920_80 vdd_M3_3920_160 3.2
c766 vdd_M3_3920_80 0 0.008f
c767 vdd_M3_3920_160 0 0.008f
r414 vdd_M3_3920_160 vdd_M3_3920_168 0.32
c768 vdd_M3_3920_160 0 0.0008f
c769 vdd_M3_3920_168 0 0.0008f
r415 vdd_M3_3920_168 vdd_M3_3920_248 3.2
c770 vdd_M3_3920_168 0 0.008f
c771 vdd_M3_3920_248 0 0.008f
r416 vdd_M3_3920_248 vdd_M3_3920_328 3.2
c772 vdd_M3_3920_248 0 0.008f
c773 vdd_M3_3920_328 0 0.008f
r417 vdd_M3_3920_328 vdd_M3_3920_336 0.32
c774 vdd_M3_3920_328 0 0.0008f
c775 vdd_M3_3920_336 0 0.0008f
r418 vdd_M3_3920_336 vdd_M3_3920_372 1.44
c776 vdd_M3_3920_336 0 0.0036f
c777 vdd_M3_3920_372 0 0.0036f
r419 vdd_M3_3760_132 vdd_M3_3760_168 1.44
c778 vdd_M3_3760_132 0 0.0036f
c779 vdd_M3_3760_168 0 0.0036f
r420 vdd_M3_3760_168 vdd_M3_3760_248 3.2
c780 vdd_M3_3760_168 0 0.008f
c781 vdd_M3_3760_248 0 0.008f
r421 vdd_M3_3760_248 vdd_M3_3760_328 3.2
c782 vdd_M3_3760_248 0 0.008f
c783 vdd_M3_3760_328 0 0.008f
r422 vdd_M3_3760_328 vdd_M3_3760_336 0.32
c784 vdd_M3_3760_328 0 0.0008f
c785 vdd_M3_3760_336 0 0.0008f
r423 vdd_M3_3760_336 vdd_M3_3760_416 3.2
c786 vdd_M3_3760_336 0 0.008f
c787 vdd_M3_3760_416 0 0.008f
r424 vdd_M3_3760_416 vdd_M3_3760_441 1.0
c788 vdd_M3_3760_416 0 0.0025000000000000005f
c789 vdd_M3_3760_441 0 0.0025000000000000005f
r425 net8_M3_3840_216 net8_M3_3840_252 1.44
c790 net8_M3_3840_216 0 0.0036f
c791 net8_M3_3840_252 0 0.0036f
r426 net8_M3_3840_252 net8_M3_3840_332 3.2
c792 net8_M3_3840_252 0 0.008f
c793 net8_M3_3840_332 0 0.008f
r427 net8_M3_3840_332 net8_M3_3840_412 3.2
c794 net8_M3_3840_332 0 0.008f
c795 net8_M3_3840_412 0 0.008f
r428 net8_M3_3840_412 net8_M3_3840_420 0.32
c796 net8_M3_3840_412 0 0.0008f
c797 net8_M3_3840_420 0 0.0008f
r429 net8_M3_3840_420 net8_M3_3840_456 1.44
c798 net8_M3_3840_420 0 0.0036f
c799 net8_M3_3840_456 0 0.0036f
r430 net8_M3_3680_216 net8_M3_3680_252 1.44
c800 net8_M3_3680_216 0 0.0036f
c801 net8_M3_3680_252 0 0.0036f
r431 net8_M3_3680_252 net8_M3_3680_332 3.2
c802 net8_M3_3680_252 0 0.008f
c803 net8_M3_3680_332 0 0.008f
r432 net8_M3_3680_332 net8_M3_3680_412 3.2
c804 net8_M3_3680_332 0 0.008f
c805 net8_M3_3680_412 0 0.008f
r433 net8_M3_3680_412 net8_M3_3680_420 0.32
c806 net8_M3_3680_412 0 0.0008f
c807 net8_M3_3680_420 0 0.0008f
r434 net8_M3_3680_420 net8_M3_3680_500 3.2
c808 net8_M3_3680_420 0 0.008f
c809 net8_M3_3680_500 0 0.008f
r435 net8_M3_3680_500 net8_M3_3680_525 1.0
c810 net8_M3_3680_500 0 0.0025000000000000005f
c811 net8_M3_3680_525 0 0.0025000000000000005f
r436 vdd_M3_3280_132 vdd_M3_3280_168 1.44
c812 vdd_M3_3280_132 0 0.0036f
c813 vdd_M3_3280_168 0 0.0036f
r437 vdd_M3_3280_168 vdd_M3_3280_248 3.2
c814 vdd_M3_3280_168 0 0.008f
c815 vdd_M3_3280_248 0 0.008f
r438 vdd_M3_3280_248 vdd_M3_3280_328 3.2
c816 vdd_M3_3280_248 0 0.008f
c817 vdd_M3_3280_328 0 0.008f
r439 vdd_M3_3280_328 vdd_M3_3280_408 3.2
c818 vdd_M3_3280_328 0 0.008f
c819 vdd_M3_3280_408 0 0.008f
r440 vdd_M3_3280_408 vdd_M3_3280_420 0.48
c820 vdd_M3_3280_408 0 0.0012000000000000001f
c821 vdd_M3_3280_420 0 0.0012000000000000001f
r441 vdd_M3_3280_420 vdd_M3_3280_456 1.44
c822 vdd_M3_3280_420 0 0.0036f
c823 vdd_M3_3280_456 0 0.0036f
r442 vdd_M3_3040_132 vdd_M3_3040_168 1.44
c824 vdd_M3_3040_132 0 0.0036f
c825 vdd_M3_3040_168 0 0.0036f
r443 vdd_M3_3040_168 vdd_M3_3040_248 3.2
c826 vdd_M3_3040_168 0 0.008f
c827 vdd_M3_3040_248 0 0.008f
r444 vdd_M3_3040_248 vdd_M3_3040_328 3.2
c828 vdd_M3_3040_248 0 0.008f
c829 vdd_M3_3040_328 0 0.008f
r445 vdd_M3_3040_328 vdd_M3_3040_336 0.32
c830 vdd_M3_3040_328 0 0.0008f
c831 vdd_M3_3040_336 0 0.0008f
r446 vdd_M3_3040_336 vdd_M3_3040_416 3.2
c832 vdd_M3_3040_336 0 0.008f
c833 vdd_M3_3040_416 0 0.008f
r447 vdd_M3_3040_416 vdd_M3_3040_420 0.16
c834 vdd_M3_3040_416 0 0.0004f
c835 vdd_M3_3040_420 0 0.0004f
r448 vdd_M3_3040_420 vdd_M3_3040_456 1.44
c836 vdd_M3_3040_420 0 0.0036f
c837 vdd_M3_3040_456 0 0.0036f
r449 vout_M3_3200_216 vout_M3_3200_252 1.44
c838 vout_M3_3200_216 0 0.0036f
c839 vout_M3_3200_252 0 0.0036f
r450 vout_M3_3200_252 vout_M3_3200_332 3.2
c840 vout_M3_3200_252 0 0.008f
c841 vout_M3_3200_332 0 0.008f
r451 vout_M3_3200_332 vout_M3_3200_412 3.2
c842 vout_M3_3200_332 0 0.008f
c843 vout_M3_3200_412 0 0.008f
r452 vout_M3_3200_412 vout_M3_3200_492 3.2
c844 vout_M3_3200_412 0 0.008f
c845 vout_M3_3200_492 0 0.008f
r453 vout_M3_3200_492 vout_M3_3200_504 0.48
c846 vout_M3_3200_492 0 0.0012000000000000001f
c847 vout_M3_3200_504 0 0.0012000000000000001f
r454 vout_M3_3200_504 vout_M3_3200_540 1.44
c848 vout_M3_3200_504 0 0.0036f
c849 vout_M3_3200_540 0 0.0036f
r455 vout_M3_2960_48 vout_M3_2960_84 1.44
c850 vout_M3_2960_48 0 0.0036f
c851 vout_M3_2960_84 0 0.0036f
r456 vout_M3_2960_84 vout_M3_2960_164 3.2
c852 vout_M3_2960_84 0 0.008f
c853 vout_M3_2960_164 0 0.008f
r457 vout_M3_2960_164 vout_M3_2960_244 3.2
c854 vout_M3_2960_164 0 0.008f
c855 vout_M3_2960_244 0 0.008f
r458 vout_M3_2960_244 vout_M3_2960_252 0.32
c856 vout_M3_2960_244 0 0.0008f
c857 vout_M3_2960_252 0 0.0008f
r459 vout_M3_2960_252 vout_M3_2960_332 3.2
c858 vout_M3_2960_252 0 0.008f
c859 vout_M3_2960_332 0 0.008f
r460 vout_M3_2960_332 vout_M3_2960_412 3.2
c860 vout_M3_2960_332 0 0.008f
c861 vout_M3_2960_412 0 0.008f
r461 vout_M3_2960_412 vout_M3_2960_492 3.2
c862 vout_M3_2960_412 0 0.008f
c863 vout_M3_2960_492 0 0.008f
r462 vout_M3_2960_492 vout_M3_2960_504 0.48
c864 vout_M3_2960_492 0 0.0012000000000000001f
c865 vout_M3_2960_504 0 0.0012000000000000001f
r463 vout_M3_2960_504 vout_M3_2960_540 1.44
c866 vout_M3_2960_504 0 0.0036f
c867 vout_M3_2960_540 0 0.0036f
r464 net8_M3_3120_300 net8_M3_3120_336 1.44
c868 net8_M3_3120_300 0 0.0036f
c869 net8_M3_3120_336 0 0.0036f
r465 net8_M3_3120_336 net8_M3_3120_416 3.2
c870 net8_M3_3120_336 0 0.008f
c871 net8_M3_3120_416 0 0.008f
r466 net8_M3_3120_416 net8_M3_3120_496 3.2
c872 net8_M3_3120_416 0 0.008f
c873 net8_M3_3120_496 0 0.008f
r467 net8_M3_3120_496 net8_M3_3120_576 3.2
c874 net8_M3_3120_496 0 0.008f
c875 net8_M3_3120_576 0 0.008f
r468 net8_M3_3120_576 net8_M3_3120_588 0.48
c876 net8_M3_3120_576 0 0.0012000000000000001f
c877 net8_M3_3120_588 0 0.0012000000000000001f
r469 net8_M3_3120_588 net8_M3_3120_624 1.44
c878 net8_M3_3120_588 0 0.0036f
c879 net8_M3_3120_624 0 0.0036f
r470 net8_M3_2880_300 net8_M3_2880_336 1.44
c880 net8_M3_2880_300 0 0.0036f
c881 net8_M3_2880_336 0 0.0036f
r471 net8_M3_2880_336 net8_M3_2880_416 3.2
c882 net8_M3_2880_336 0 0.008f
c883 net8_M3_2880_416 0 0.008f
r472 net8_M3_2880_416 net8_M3_2880_420 0.16
c884 net8_M3_2880_416 0 0.0004f
c885 net8_M3_2880_420 0 0.0004f
r473 net8_M3_2880_420 net8_M3_2880_500 3.2
c886 net8_M3_2880_420 0 0.008f
c887 net8_M3_2880_500 0 0.008f
r474 net8_M3_2880_500 net8_M3_2880_504 0.16
c888 net8_M3_2880_500 0 0.0004f
c889 net8_M3_2880_504 0 0.0004f
r475 net8_M3_2880_504 net8_M3_2880_584 3.2
c890 net8_M3_2880_504 0 0.008f
c891 net8_M3_2880_584 0 0.008f
r476 net8_M3_2880_584 net8_M3_2880_588 0.16
c892 net8_M3_2880_584 0 0.0004f
c893 net8_M3_2880_588 0 0.0004f
r477 net8_M3_2880_588 net8_M3_2880_624 1.44
c894 net8_M3_2880_588 0 0.0036f
c895 net8_M3_2880_624 0 0.0036f
r478 vss_M3_560_132 vss_M3_560_168 1.44
c896 vss_M3_560_132 0 0.0036f
c897 vss_M3_560_168 0 0.0036f
r479 vss_M3_560_168 vss_M3_560_248 3.2
c898 vss_M3_560_168 0 0.008f
c899 vss_M3_560_248 0 0.008f
r480 vss_M3_560_248 vss_M3_560_328 3.2
c900 vss_M3_560_248 0 0.008f
c901 vss_M3_560_328 0 0.008f
r481 vss_M3_560_328 vss_M3_560_408 3.2
c902 vss_M3_560_328 0 0.008f
c903 vss_M3_560_408 0 0.008f
r482 vss_M3_560_408 vss_M3_560_420 0.48
c904 vss_M3_560_408 0 0.0012000000000000001f
c905 vss_M3_560_420 0 0.0012000000000000001f
r483 vss_M3_560_420 vss_M3_560_456 1.44
c906 vss_M3_560_420 0 0.0036f
c907 vss_M3_560_456 0 0.0036f
r484 vss_M3_800_132 vss_M3_800_168 1.44
c908 vss_M3_800_132 0 0.0036f
c909 vss_M3_800_168 0 0.0036f
r485 vss_M3_800_168 vss_M3_800_248 3.2
c910 vss_M3_800_168 0 0.008f
c911 vss_M3_800_248 0 0.008f
r486 vss_M3_800_248 vss_M3_800_328 3.2
c912 vss_M3_800_248 0 0.008f
c913 vss_M3_800_328 0 0.008f
r487 vss_M3_800_328 vss_M3_800_408 3.2
c914 vss_M3_800_328 0 0.008f
c915 vss_M3_800_408 0 0.008f
r488 vss_M3_800_408 vss_M3_800_420 0.48
c916 vss_M3_800_408 0 0.0012000000000000001f
c917 vss_M3_800_420 0 0.0012000000000000001f
r489 vss_M3_800_420 vss_M3_800_456 1.44
c918 vss_M3_800_420 0 0.0036f
c919 vss_M3_800_456 0 0.0036f
r490 id_M3_640__36 id_M3_640_0 1.44
c920 id_M3_640__36 0 0.0036f
c921 id_M3_640_0 0 0.0036f
r491 id_M3_640_0 id_M3_640_80 3.2
c922 id_M3_640_0 0 0.008f
c923 id_M3_640_80 0 0.008f
r492 id_M3_640_80 id_M3_640_160 3.2
c924 id_M3_640_80 0 0.008f
c925 id_M3_640_160 0 0.008f
r493 id_M3_640_160 id_M3_640_240 3.2
c926 id_M3_640_160 0 0.008f
c927 id_M3_640_240 0 0.008f
r494 id_M3_640_240 id_M3_640_252 0.48
c928 id_M3_640_240 0 0.0012000000000000001f
c929 id_M3_640_252 0 0.0012000000000000001f
r495 id_M3_640_252 id_M3_640_332 3.2
c930 id_M3_640_252 0 0.008f
c931 id_M3_640_332 0 0.008f
r496 id_M3_640_332 id_M3_640_412 3.2
c932 id_M3_640_332 0 0.008f
c933 id_M3_640_412 0 0.008f
r497 id_M3_640_412 id_M3_640_492 3.2
c934 id_M3_640_412 0 0.008f
c935 id_M3_640_492 0 0.008f
r498 id_M3_640_492 id_M3_640_504 0.48
c936 id_M3_640_492 0 0.0012000000000000001f
c937 id_M3_640_504 0 0.0012000000000000001f
r499 id_M3_640_504 id_M3_640_540 1.44
c938 id_M3_640_504 0 0.0036f
c939 id_M3_640_540 0 0.0036f
r500 id_M3_880_216 id_M3_880_252 1.44
c940 id_M3_880_216 0 0.0036f
c941 id_M3_880_252 0 0.0036f
r501 id_M3_880_252 id_M3_880_332 3.2
c942 id_M3_880_252 0 0.008f
c943 id_M3_880_332 0 0.008f
r502 id_M3_880_332 id_M3_880_412 3.2
c944 id_M3_880_332 0 0.008f
c945 id_M3_880_412 0 0.008f
r503 id_M3_880_412 id_M3_880_492 3.2
c946 id_M3_880_412 0 0.008f
c947 id_M3_880_492 0 0.008f
r504 id_M3_880_492 id_M3_880_504 0.48
c948 id_M3_880_492 0 0.0012000000000000001f
c949 id_M3_880_504 0 0.0012000000000000001f
r505 id_M3_880_504 id_M3_880_540 1.44
c950 id_M3_880_504 0 0.0036f
c951 id_M3_880_540 0 0.0036f
r506 net10_M3_720_300 net10_M3_720_336 1.44
c952 net10_M3_720_300 0 0.0036f
c953 net10_M3_720_336 0 0.0036f
r507 net10_M3_720_336 net10_M3_720_416 3.2
c954 net10_M3_720_336 0 0.008f
c955 net10_M3_720_416 0 0.008f
r508 net10_M3_720_416 net10_M3_720_496 3.2
c956 net10_M3_720_416 0 0.008f
c957 net10_M3_720_496 0 0.008f
r509 net10_M3_720_496 net10_M3_720_576 3.2
c958 net10_M3_720_496 0 0.008f
c959 net10_M3_720_576 0 0.008f
r510 net10_M3_720_576 net10_M3_720_588 0.48
c960 net10_M3_720_576 0 0.0012000000000000001f
c961 net10_M3_720_588 0 0.0012000000000000001f
r511 net10_M3_720_588 net10_M3_720_624 1.44
c962 net10_M3_720_588 0 0.0036f
c963 net10_M3_720_624 0 0.0036f
r512 net10_M3_960_128 net10_M3_960_168 1.6
c964 net10_M3_960_128 0 0.004f
c965 net10_M3_960_168 0 0.004f
r513 net10_M3_960_168 net10_M3_960_248 3.2
c966 net10_M3_960_168 0 0.008f
c967 net10_M3_960_248 0 0.008f
r514 net10_M3_960_248 net10_M3_960_328 3.2
c968 net10_M3_960_248 0 0.008f
c969 net10_M3_960_328 0 0.008f
r515 net10_M3_960_328 net10_M3_960_336 0.32
c970 net10_M3_960_328 0 0.0008f
c971 net10_M3_960_336 0 0.0008f
r516 net10_M3_960_336 net10_M3_960_416 3.2
c972 net10_M3_960_336 0 0.008f
c973 net10_M3_960_416 0 0.008f
r517 net10_M3_960_416 net10_M3_960_496 3.2
c974 net10_M3_960_416 0 0.008f
c975 net10_M3_960_496 0 0.008f
r518 net10_M3_960_496 net10_M3_960_576 3.2
c976 net10_M3_960_496 0 0.008f
c977 net10_M3_960_576 0 0.008f
r519 net10_M3_960_576 net10_M3_960_588 0.48
c978 net10_M3_960_576 0 0.0012000000000000001f
c979 net10_M3_960_588 0 0.0012000000000000001f
r520 net10_M3_960_588 net10_M3_960_624 1.44
c980 net10_M3_960_588 0 0.0036f
c981 net10_M3_960_624 0 0.0036f
r521 net8_M3_2160_216 net8_M3_2160_252 1.44
c982 net8_M3_2160_216 0 0.0036f
c983 net8_M3_2160_252 0 0.0036f
r522 net8_M3_2160_252 net8_M3_2160_332 3.2
c984 net8_M3_2160_252 0 0.008f
c985 net8_M3_2160_332 0 0.008f
r523 net8_M3_2160_332 net8_M3_2160_412 3.2
c986 net8_M3_2160_332 0 0.008f
c987 net8_M3_2160_412 0 0.008f
r524 net8_M3_2160_412 net8_M3_2160_492 3.2
c988 net8_M3_2160_412 0 0.008f
c989 net8_M3_2160_492 0 0.008f
r525 net8_M3_2160_492 net8_M3_2160_504 0.48
c990 net8_M3_2160_492 0 0.0012000000000000001f
c991 net8_M3_2160_504 0 0.0012000000000000001f
r526 net8_M3_2160_504 net8_M3_2160_544 1.6
c992 net8_M3_2160_504 0 0.004f
c993 net8_M3_2160_544 0 0.004f
r527 vdd_M3_3600_231 vdd_M3_3600_311 3.2
c994 vdd_M3_3600_231 0 0.008f
c995 vdd_M3_3600_311 0 0.008f
r528 vdd_M3_3600_311 vdd_M3_3600_336 1.0
c996 vdd_M3_3600_311 0 0.0025000000000000005f
c997 vdd_M3_3600_336 0 0.0025000000000000005f
r529 vdd_M3_3600_336 vdd_M3_3600_416 3.2
c998 vdd_M3_3600_336 0 0.008f
c999 vdd_M3_3600_416 0 0.008f
r530 vdd_M3_3600_416 vdd_M3_3600_441 1.0
c1000 vdd_M3_3600_416 0 0.0025000000000000005f
c1001 vdd_M3_3600_441 0 0.0025000000000000005f
r531 vdd_M3_3360_231 vdd_M3_3360_311 3.2
c1002 vdd_M3_3360_231 0 0.008f
c1003 vdd_M3_3360_311 0 0.008f
r532 vdd_M3_3360_311 vdd_M3_3360_336 1.0
c1004 vdd_M3_3360_311 0 0.0025000000000000005f
c1005 vdd_M3_3360_336 0 0.0025000000000000005f
r533 vdd_M3_3360_336 vdd_M3_3360_416 3.2
c1006 vdd_M3_3360_336 0 0.008f
c1007 vdd_M3_3360_416 0 0.008f
r534 vdd_M3_3360_416 vdd_M3_3360_441 1.0
c1008 vdd_M3_3360_416 0 0.0025000000000000005f
c1009 vdd_M3_3360_441 0 0.0025000000000000005f
r535 vout_M3_2480_48 vout_M3_2480_84 1.44
c1010 vout_M3_2480_48 0 0.0036f
c1011 vout_M3_2480_84 0 0.0036f
r536 vout_M3_2480_84 vout_M3_2480_164 3.2
c1012 vout_M3_2480_84 0 0.008f
c1013 vout_M3_2480_164 0 0.008f
r537 vout_M3_2480_164 vout_M3_2480_244 3.2
c1014 vout_M3_2480_164 0 0.008f
c1015 vout_M3_2480_244 0 0.008f
r538 vout_M3_2480_244 vout_M3_2480_252 0.32
c1016 vout_M3_2480_244 0 0.0008f
c1017 vout_M3_2480_252 0 0.0008f
r539 vout_M3_2480_252 vout_M3_2480_332 3.2
c1018 vout_M3_2480_252 0 0.008f
c1019 vout_M3_2480_332 0 0.008f
r540 vout_M3_2480_332 vout_M3_2480_336 0.16
c1020 vout_M3_2480_332 0 0.0004f
c1021 vout_M3_2480_336 0 0.0004f
r541 vout_M3_2480_336 vout_M3_2480_372 1.44
c1022 vout_M3_2480_336 0 0.0036f
c1023 vout_M3_2480_372 0 0.0036f
r542 vout_M3_2640_147 vout_M3_2640_227 3.2
c1024 vout_M3_2640_147 0 0.008f
c1025 vout_M3_2640_227 0 0.008f
r543 vout_M3_2640_227 vout_M3_2640_252 1.0
c1026 vout_M3_2640_227 0 0.0025000000000000005f
c1027 vout_M3_2640_252 0 0.0025000000000000005f
r544 vout_M3_2640_252 vout_M3_2640_332 3.2
c1028 vout_M3_2640_252 0 0.008f
c1029 vout_M3_2640_332 0 0.008f
r545 vout_M3_2640_332 vout_M3_2640_357 1.0
c1030 vout_M3_2640_332 0 0.0025000000000000005f
c1031 vout_M3_2640_357 0 0.0025000000000000005f
r546 vout_M3_2400__36 vout_M3_2400_0 1.44
c1032 vout_M3_2400__36 0 0.0036f
c1033 vout_M3_2400_0 0 0.0036f
r547 vout_M3_2400_0 vout_M3_2400_80 3.2
c1034 vout_M3_2400_0 0 0.008f
c1035 vout_M3_2400_80 0 0.008f
r548 vout_M3_2400_80 vout_M3_2400_160 3.2
c1036 vout_M3_2400_80 0 0.008f
c1037 vout_M3_2400_160 0 0.008f
r549 vout_M3_2400_160 vout_M3_2400_240 3.2
c1038 vout_M3_2400_160 0 0.008f
c1039 vout_M3_2400_240 0 0.008f
r550 vout_M3_2400_240 vout_M3_2400_252 0.48
c1040 vout_M3_2400_240 0 0.0012000000000000001f
c1041 vout_M3_2400_252 0 0.0012000000000000001f
r551 vout_M3_2400_252 vout_M3_2400_288 1.44
c1042 vout_M3_2400_252 0 0.0036f
c1043 vout_M3_2400_288 0 0.0036f
r552 net10_M3_1280_63 net10_M3_1280_143 3.2
c1044 net10_M3_1280_63 0 0.008f
c1045 net10_M3_1280_143 0 0.008f
r553 net10_M3_1280_143 net10_M3_1280_168 1.0
c1046 net10_M3_1280_143 0 0.0025000000000000005f
c1047 net10_M3_1280_168 0 0.0025000000000000005f
r554 net10_M3_1280_168 net10_M3_1280_248 3.2
c1048 net10_M3_1280_168 0 0.008f
c1049 net10_M3_1280_248 0 0.008f
r555 net10_M3_1280_248 net10_M3_1280_273 1.0
c1050 net10_M3_1280_248 0 0.0025000000000000005f
c1051 net10_M3_1280_273 0 0.0025000000000000005f
r556 vinp_M3_1920_128 vinp_M3_1920_168 1.6
c1052 vinp_M3_1920_128 0 0.004f
c1053 vinp_M3_1920_168 0 0.004f
r557 vinp_M3_1920_168 vinp_M3_1920_248 3.2
c1054 vinp_M3_1920_168 0 0.008f
c1055 vinp_M3_1920_248 0 0.008f
r558 vinp_M3_1920_248 vinp_M3_1920_328 3.2
c1056 vinp_M3_1920_248 0 0.008f
c1057 vinp_M3_1920_328 0 0.008f
r559 vinp_M3_1920_328 vinp_M3_1920_408 3.2
c1058 vinp_M3_1920_328 0 0.008f
c1059 vinp_M3_1920_408 0 0.008f
r560 vinp_M3_1920_408 vinp_M3_1920_420 0.48
c1060 vinp_M3_1920_408 0 0.0012000000000000001f
c1061 vinp_M3_1920_420 0 0.0012000000000000001f
r561 vinp_M3_1920_420 vinp_M3_1920_456 1.44
c1062 vinp_M3_1920_420 0 0.0036f
c1063 vinp_M3_1920_456 0 0.0036f
r562 vinp_M3_1600__40 vinp_M3_1600_0 1.6
c1064 vinp_M3_1600__40 0 0.004f
c1065 vinp_M3_1600_0 0 0.004f
r563 vinp_M3_1600_0 vinp_M3_1600_80 3.2
c1066 vinp_M3_1600_0 0 0.008f
c1067 vinp_M3_1600_80 0 0.008f
r564 vinp_M3_1600_80 vinp_M3_1600_160 3.2
c1068 vinp_M3_1600_80 0 0.008f
c1069 vinp_M3_1600_160 0 0.008f
r565 vinp_M3_1600_160 vinp_M3_1600_240 3.2
c1070 vinp_M3_1600_160 0 0.008f
c1071 vinp_M3_1600_240 0 0.008f
r566 vinp_M3_1600_240 vinp_M3_1600_252 0.48
c1072 vinp_M3_1600_240 0 0.0012000000000000001f
c1073 vinp_M3_1600_252 0 0.0012000000000000001f
r567 vinp_M3_1600_252 vinp_M3_1600_288 1.44
c1074 vinp_M3_1600_252 0 0.0036f
c1075 vinp_M3_1600_288 0 0.0036f
r568 vinp_M3_1360__36 vinp_M3_1360_0 1.44
c1076 vinp_M3_1360__36 0 0.0036f
c1077 vinp_M3_1360_0 0 0.0036f
r569 vinp_M3_1360_0 vinp_M3_1360_80 3.2
c1078 vinp_M3_1360_0 0 0.008f
c1079 vinp_M3_1360_80 0 0.008f
r570 vinp_M3_1360_80 vinp_M3_1360_160 3.2
c1080 vinp_M3_1360_80 0 0.008f
c1081 vinp_M3_1360_160 0 0.008f
r571 vinp_M3_1360_160 vinp_M3_1360_240 3.2
c1082 vinp_M3_1360_160 0 0.008f
c1083 vinp_M3_1360_240 0 0.008f
r572 vinp_M3_1360_240 vinp_M3_1360_252 0.48
c1084 vinp_M3_1360_240 0 0.0012000000000000001f
c1085 vinp_M3_1360_252 0 0.0012000000000000001f
r573 vinp_M3_1360_252 vinp_M3_1360_288 1.44
c1086 vinp_M3_1360_252 0 0.0036f
c1087 vinp_M3_1360_288 0 0.0036f
r574 vdd_M2_3920_0 vdd_M3_3920_0 50
r575 vdd_M2_3920_168 vdd_M3_3920_168 50
r576 vdd_M2_3920_336 vdd_M3_3920_336 50
r577 vdd_M2_3760_168 vdd_M3_3760_168 50
r578 vdd_M2_3760_336 vdd_M3_3760_336 50
r579 net8_M2_3840_252 net8_M3_3840_252 50
r580 net8_M2_3840_420 net8_M3_3840_420 50
r581 net8_M2_3680_252 net8_M3_3680_252 50
r582 net8_M2_3680_420 net8_M3_3680_420 50
r583 vdd_M2_3280_168 vdd_M3_3280_168 50
r584 vdd_M2_3280_420 vdd_M3_3280_420 50
r585 vdd_M2_3040_168 vdd_M3_3040_168 50
r586 vdd_M2_3040_420 vdd_M3_3040_420 50
r587 vout_M2_3200_252 vout_M3_3200_252 50
r588 vout_M2_3200_504 vout_M3_3200_504 50
r589 vout_M2_2960_84 vout_M3_2960_84 50
r590 vout_M2_2960_252 vout_M3_2960_252 50
r591 vout_M2_2960_504 vout_M3_2960_504 50
r592 net8_M2_3120_336 net8_M3_3120_336 50
r593 net8_M2_3120_588 net8_M3_3120_588 50
r594 net8_M2_2880_336 net8_M3_2880_336 50
r595 net8_M2_2880_588 net8_M3_2880_588 50
r596 vss_M2_560_168 vss_M3_560_168 50
r597 vss_M2_560_420 vss_M3_560_420 50
r598 vss_M2_800_168 vss_M3_800_168 50
r599 vss_M2_800_420 vss_M3_800_420 50
r600 id_M2_640_0 id_M3_640_0 50
r601 id_M2_640_252 id_M3_640_252 50
r602 id_M2_640_504 id_M3_640_504 50
r603 id_M2_880_252 id_M3_880_252 50
r604 id_M2_880_504 id_M3_880_504 50
r605 net10_M2_720_336 net10_M3_720_336 50
r606 net10_M2_720_588 net10_M3_720_588 50
r607 net10_M2_960_336 net10_M3_960_336 50
r608 net10_M2_960_588 net10_M3_960_588 50
r609 net8_M2_2160_252 net8_M3_2160_252 50
r610 vdd_M2_3360_336 vdd_M3_3360_336 50
r611 vdd_M2_3600_336 vdd_M3_3600_336 50
r612 vout_M2_2400_0 vout_M3_2400_0 50
r613 vout_M2_2400_252 vout_M3_2400_252 50
r614 vout_M2_2480_84 vout_M3_2480_84 50
r615 vout_M2_2480_336 vout_M3_2480_336 50
r616 vout_M2_2640_252 vout_M3_2640_252 50
r617 net10_M2_1280_168 net10_M3_1280_168 50
r618 vinp_M2_1360_0 vinp_M3_1360_0 50
r619 vinp_M2_1360_252 vinp_M3_1360_252 50
r620 vinp_M2_1600_252 vinp_M3_1600_252 50
r621 vinp_M2_1920_420 vinp_M3_1920_420 50
r622 net8_M4_2840_420 net8_M4_2880_420 1.2
c1088 net8_M4_2840_420 0 0.004f
c1089 net8_M4_2880_420 0 0.004f
r623 net8_M4_2880_420 net8_M4_2960_420 2.4
c1090 net8_M4_2880_420 0 0.008f
c1091 net8_M4_2960_420 0 0.008f
r624 net8_M4_2960_420 net8_M4_3040_420 2.4
c1092 net8_M4_2960_420 0 0.008f
c1093 net8_M4_3040_420 0 0.008f
r625 net8_M4_3040_420 net8_M4_3120_420 2.4
c1094 net8_M4_3040_420 0 0.008f
c1095 net8_M4_3120_420 0 0.008f
r626 net8_M4_3120_420 net8_M4_3200_420 2.4
c1096 net8_M4_3120_420 0 0.008f
c1097 net8_M4_3200_420 0 0.008f
r627 net8_M4_3200_420 net8_M4_3280_420 2.4
c1098 net8_M4_3200_420 0 0.008f
c1099 net8_M4_3280_420 0 0.008f
r628 net8_M4_3280_420 net8_M4_3360_420 2.4
c1100 net8_M4_3280_420 0 0.008f
c1101 net8_M4_3360_420 0 0.008f
r629 net8_M4_3360_420 net8_M4_3440_420 2.4
c1102 net8_M4_3360_420 0 0.008f
c1103 net8_M4_3440_420 0 0.008f
r630 net8_M4_3440_420 net8_M4_3520_420 2.4
c1104 net8_M4_3440_420 0 0.008f
c1105 net8_M4_3520_420 0 0.008f
r631 net8_M4_3520_420 net8_M4_3600_420 2.4
c1106 net8_M4_3520_420 0 0.008f
c1107 net8_M4_3600_420 0 0.008f
r632 net8_M4_3600_420 net8_M4_3680_420 2.4
c1108 net8_M4_3600_420 0 0.008f
c1109 net8_M4_3680_420 0 0.008f
r633 net8_M4_3680_420 net8_M4_3720_420 1.2
c1110 net8_M4_3680_420 0 0.004f
c1111 net8_M4_3720_420 0 0.004f
r634 net8_M4_2120_504 net8_M4_2160_504 1.2
c1112 net8_M4_2120_504 0 0.004f
c1113 net8_M4_2160_504 0 0.004f
r635 net8_M4_2160_504 net8_M4_2240_504 2.4
c1114 net8_M4_2160_504 0 0.008f
c1115 net8_M4_2240_504 0 0.008f
r636 net8_M4_2240_504 net8_M4_2320_504 2.4
c1116 net8_M4_2240_504 0 0.008f
c1117 net8_M4_2320_504 0 0.008f
r637 net8_M4_2320_504 net8_M4_2400_504 2.4
c1118 net8_M4_2320_504 0 0.008f
c1119 net8_M4_2400_504 0 0.008f
r638 net8_M4_2400_504 net8_M4_2480_504 2.4
c1120 net8_M4_2400_504 0 0.008f
c1121 net8_M4_2480_504 0 0.008f
r639 net8_M4_2480_504 net8_M4_2560_504 2.4
c1122 net8_M4_2480_504 0 0.008f
c1123 net8_M4_2560_504 0 0.008f
r640 net8_M4_2560_504 net8_M4_2640_504 2.4
c1124 net8_M4_2560_504 0 0.008f
c1125 net8_M4_2640_504 0 0.008f
r641 net8_M4_2640_504 net8_M4_2720_504 2.4
c1126 net8_M4_2640_504 0 0.008f
c1127 net8_M4_2720_504 0 0.008f
r642 net8_M4_2720_504 net8_M4_2800_504 2.4
c1128 net8_M4_2720_504 0 0.008f
c1129 net8_M4_2800_504 0 0.008f
r643 net8_M4_2800_504 net8_M4_2880_504 2.4
c1130 net8_M4_2800_504 0 0.008f
c1131 net8_M4_2880_504 0 0.008f
r644 net8_M4_2880_504 net8_M4_2920_504 1.2
c1132 net8_M4_2880_504 0 0.004f
c1133 net8_M4_2920_504 0 0.004f
r645 vdd_M4_3000_336 vdd_M4_3040_336 1.2
c1134 vdd_M4_3000_336 0 0.004f
c1135 vdd_M4_3040_336 0 0.004f
r646 vdd_M4_3040_336 vdd_M4_3120_336 2.4
c1136 vdd_M4_3040_336 0 0.008f
c1137 vdd_M4_3120_336 0 0.008f
r647 vdd_M4_3120_336 vdd_M4_3200_336 2.4
c1138 vdd_M4_3120_336 0 0.008f
c1139 vdd_M4_3200_336 0 0.008f
r648 vdd_M4_3200_336 vdd_M4_3280_336 2.4
c1140 vdd_M4_3200_336 0 0.008f
c1141 vdd_M4_3280_336 0 0.008f
r649 vdd_M4_3280_336 vdd_M4_3360_336 2.4
c1142 vdd_M4_3280_336 0 0.008f
c1143 vdd_M4_3360_336 0 0.008f
r650 vdd_M4_3360_336 vdd_M4_3400_336 1.2
c1144 vdd_M4_3360_336 0 0.004f
c1145 vdd_M4_3400_336 0 0.004f
r651 vdd_M4_3560_336 vdd_M4_3600_336 1.2
c1146 vdd_M4_3560_336 0 0.004f
c1147 vdd_M4_3600_336 0 0.004f
r652 vdd_M4_3600_336 vdd_M4_3680_336 2.4
c1148 vdd_M4_3600_336 0 0.008f
c1149 vdd_M4_3680_336 0 0.008f
r653 vdd_M4_3680_336 vdd_M4_3760_336 2.4
c1150 vdd_M4_3680_336 0 0.008f
c1151 vdd_M4_3760_336 0 0.008f
r654 vdd_M4_3760_336 vdd_M4_3800_336 1.2
c1152 vdd_M4_3760_336 0 0.004f
c1153 vdd_M4_3800_336 0 0.004f
r655 vout_M4_2440_252 vout_M4_2480_252 1.2
c1154 vout_M4_2440_252 0 0.004f
c1155 vout_M4_2480_252 0 0.004f
r656 vout_M4_2480_252 vout_M4_2560_252 2.4
c1156 vout_M4_2480_252 0 0.008f
c1157 vout_M4_2560_252 0 0.008f
r657 vout_M4_2560_252 vout_M4_2640_252 2.4
c1158 vout_M4_2560_252 0 0.008f
c1159 vout_M4_2640_252 0 0.008f
r658 vout_M4_2640_252 vout_M4_2680_252 1.2
c1160 vout_M4_2640_252 0 0.004f
c1161 vout_M4_2680_252 0 0.004f
r659 net10_M4_920_168 net10_M4_960_168 1.2
c1162 net10_M4_920_168 0 0.004f
c1163 net10_M4_960_168 0 0.004f
r660 net10_M4_960_168 net10_M4_1040_168 2.4
c1164 net10_M4_960_168 0 0.008f
c1165 net10_M4_1040_168 0 0.008f
r661 net10_M4_1040_168 net10_M4_1120_168 2.4
c1166 net10_M4_1040_168 0 0.008f
c1167 net10_M4_1120_168 0 0.008f
r662 net10_M4_1120_168 net10_M4_1200_168 2.4
c1168 net10_M4_1120_168 0 0.008f
c1169 net10_M4_1200_168 0 0.008f
r663 net10_M4_1200_168 net10_M4_1280_168 2.4
c1170 net10_M4_1200_168 0 0.008f
c1171 net10_M4_1280_168 0 0.008f
r664 net10_M4_1280_168 net10_M4_1320_168 1.2
c1172 net10_M4_1280_168 0 0.004f
c1173 net10_M4_1320_168 0 0.004f
r665 vinp_M4_1400_168 vinp_M4_1440_168 1.2
c1174 vinp_M4_1400_168 0 0.004f
c1175 vinp_M4_1440_168 0 0.004f
r666 vinp_M4_1440_168 vinp_M4_1520_168 2.4
c1176 vinp_M4_1440_168 0 0.008f
c1177 vinp_M4_1520_168 0 0.008f
r667 vinp_M4_1520_168 vinp_M4_1600_168 2.4
c1178 vinp_M4_1520_168 0 0.008f
c1179 vinp_M4_1600_168 0 0.008f
r668 vinp_M4_1600_168 vinp_M4_1680_168 2.4
c1180 vinp_M4_1600_168 0 0.008f
c1181 vinp_M4_1680_168 0 0.008f
r669 vinp_M4_1680_168 vinp_M4_1760_168 2.4
c1182 vinp_M4_1680_168 0 0.008f
c1183 vinp_M4_1760_168 0 0.008f
r670 vinp_M4_1760_168 vinp_M4_1840_168 2.4
c1184 vinp_M4_1760_168 0 0.008f
c1185 vinp_M4_1840_168 0 0.008f
r671 vinp_M4_1840_168 vinp_M4_1920_168 2.4
c1186 vinp_M4_1840_168 0 0.008f
c1187 vinp_M4_1920_168 0 0.008f
r672 vinp_M4_1920_168 vinp_M4_1960_168 1.2
c1188 vinp_M4_1920_168 0 0.004f
c1189 vinp_M4_1960_168 0 0.004f
r673 vinp_M4_1400_0 vinp_M4_1440_0 1.2
c1190 vinp_M4_1400_0 0 0.004f
c1191 vinp_M4_1440_0 0 0.004f
r674 vinp_M4_1440_0 vinp_M4_1520_0 2.4
c1192 vinp_M4_1440_0 0 0.008f
c1193 vinp_M4_1520_0 0 0.008f
r675 vinp_M4_1520_0 vinp_M4_1600_0 2.4
c1194 vinp_M4_1520_0 0 0.008f
c1195 vinp_M4_1600_0 0 0.008f
r676 vinp_M4_1600_0 vinp_M4_1640_0 1.2
c1196 vinp_M4_1600_0 0 0.004f
c1197 vinp_M4_1640_0 0 0.004f
r677 net8_M3_2160_504 net8_M4_2160_504 50
r678 net8_M3_2880_420 net8_M4_2880_420 50
r679 net8_M3_2880_504 net8_M4_2880_504 50
r680 net8_M3_3680_420 net8_M4_3680_420 50
r681 vdd_M3_3040_336 vdd_M4_3040_336 50
r682 vdd_M3_3360_336 vdd_M4_3360_336 50
r683 vdd_M3_3600_336 vdd_M4_3600_336 50
r684 vdd_M3_3760_336 vdd_M4_3760_336 50
r685 vout_M3_2480_252 vout_M4_2480_252 50
r686 vout_M3_2640_252 vout_M4_2640_252 50
r687 net10_M3_960_168 net10_M4_960_168 50
r688 net10_M3_1280_168 net10_M4_1280_168 50
r689 vinp_M3_1600_0 vinp_M4_1600_0 50
r690 vinp_M3_1920_168 vinp_M4_1920_168 50
r691 vinp_M5_1440__40 vinp_M5_1440_0 0.8
c1198 vinp_M5_1440__40 0 0.004f
c1199 vinp_M5_1440_0 0 0.004f
r692 vinp_M5_1440_0 vinp_M5_1440_80 1.6
c1200 vinp_M5_1440_0 0 0.008f
c1201 vinp_M5_1440_80 0 0.008f
r693 vinp_M5_1440_80 vinp_M5_1440_160 1.6
c1202 vinp_M5_1440_80 0 0.008f
c1203 vinp_M5_1440_160 0 0.008f
r694 vinp_M5_1440_160 vinp_M5_1440_168 0.16
c1204 vinp_M5_1440_160 0 0.0008f
c1205 vinp_M5_1440_168 0 0.0008f
r695 vinp_M5_1440_168 vinp_M5_1440_208 0.8
c1206 vinp_M5_1440_168 0 0.004f
c1207 vinp_M5_1440_208 0 0.004f
r696 vinp_M4_1440_0 vinp_M5_1440_0 50
r697 vinp_M4_1440_168 vinp_M5_1440_168 50
r698 net_m1_M1_X0_Y0_G net8_M1_3840_168 50
r699 net_m1_M1_X0_Y0_S vdd_M1_3920_336 50
r700 net_m1_M1_X0_Y0_S vdd_M1_3920_462 50
r701 net_m1_M1_X0_Y0_S vdd_M1_3920_588 50
r702 net_m1_M1_X0_Y0_D net8_M1_3760_336 50
r703 net_m1_M1_X0_Y0_D net8_M1_3760_462 50
r704 net_m1_M1_X0_Y0_D net8_M1_3760_588 50
r705 net_m2_M1_X0_Y0_G net8_M1_3120_168 50
r706 net_m2_M1_X0_Y0_S vdd_M1_3200_336 50
r707 net_m2_M1_X0_Y0_S vdd_M1_3200_462 50
r708 net_m2_M1_X0_Y0_S vdd_M1_3200_588 50
r709 net_m2_M1_X0_Y0_D vout_M1_3040_336 50
r710 net_m2_M1_X0_Y0_D vout_M1_3040_462 50
r711 net_m2_M1_X0_Y0_D vout_M1_3040_588 50
r712 net_m5_m4_M1_X0_Y0_G id_M1_400_168 50
r713 net_m5_m4_M1_X0_Y0_S vss_M1_320_336 50
r714 net_m5_m4_M1_X0_Y0_S vss_M1_320_462 50
r715 net_m5_m4_M1_X0_Y0_S vss_M1_320_588 50
r716 net_m5_m4_M1_X0_Y0_D id_M1_480_336 50
r717 net_m5_m4_M1_X0_Y0_D id_M1_480_462 50
r718 net_m5_m4_M1_X0_Y0_D id_M1_480_588 50
r719 net_m5_m4_M2_X1_Y0_G id_M1_1040_168 50
r720 net_m5_m4_M2_X1_Y0_S vss_M1_960_336 50
r721 net_m5_m4_M2_X1_Y0_S vss_M1_960_462 50
r722 net_m5_m4_M2_X1_Y0_S vss_M1_960_588 50
r723 net_m5_m4_M2_X1_Y0_D net10_M1_1120_336 50
r724 net_m5_m4_M2_X1_Y0_D net10_M1_1120_462 50
r725 net_m5_m4_M2_X1_Y0_D net10_M1_1120_588 50
r726 net_m0_m3_M1_X0_Y0_G vinp_M1_1760_168 50
r727 net_m0_m3_M1_X0_Y0_S net10_M1_1680_336 50
r728 net_m0_m3_M1_X0_Y0_S net10_M1_1680_462 50
r729 net_m0_m3_M1_X0_Y0_S net10_M1_1680_588 50
r730 net_m0_m3_M1_X0_Y0_D net8_M1_1840_336 50
r731 net_m0_m3_M1_X0_Y0_D net8_M1_1840_462 50
r732 net_m0_m3_M1_X0_Y0_D net8_M1_1840_588 50
r733 net_m0_m3_M2_X1_Y0_G vinn_M1_2400_168 50
r734 net_m0_m3_M2_X1_Y0_S net10_M1_2320_336 50
r735 net_m0_m3_M2_X1_Y0_S net10_M1_2320_462 50
r736 net_m0_m3_M2_X1_Y0_S net10_M1_2320_588 50
r737 net_m0_m3_M2_X1_Y0_D vout_M1_2480_336 50
r738 net_m0_m3_M2_X1_Y0_D vout_M1_2480_462 50
r739 net_m0_m3_M2_X1_Y0_D vout_M1_2480_588 50

x_m1_M1_X0_Y0_0 net_m1_M1_X0_Y0_D net_m1_M1_X0_Y0_G net_m1_M1_X0_Y0_diff vdd! pmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m1_M1_X0_Y0_1 net_m1_M1_X0_Y0_diff net_m1_M1_X0_Y0_G net_m1_M1_X0_Y0_S vdd! pmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m2_M1_X0_Y0_0 net_m2_M1_X0_Y0_D net_m2_M1_X0_Y0_G net_m2_M1_X0_Y0_diff vdd! pmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m2_M1_X0_Y0_1 net_m2_M1_X0_Y0_diff net_m2_M1_X0_Y0_G net_m2_M1_X0_Y0_S vdd! pmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m5_m4_M1_X0_Y0_0 net_m5_m4_M1_X0_Y0_D net_m5_m4_M1_X0_Y0_G net_m5_m4_M1_X0_Y0_diff gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m5_m4_M1_X0_Y0_1 net_m5_m4_M1_X0_Y0_diff net_m5_m4_M1_X0_Y0_G net_m5_m4_M1_X0_Y0_S gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m5_m4_M2_X1_Y0_0 net_m5_m4_M2_X1_Y0_D net_m5_m4_M2_X1_Y0_G net_m5_m4_M2_X1_Y0_diff gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m5_m4_M2_X1_Y0_1 net_m5_m4_M2_X1_Y0_diff net_m5_m4_M2_X1_Y0_G net_m5_m4_M2_X1_Y0_S gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m0_m3_M1_X0_Y0_0 net_m0_m3_M1_X0_Y0_D net_m0_m3_M1_X0_Y0_G net_m0_m3_M1_X0_Y0_diff gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m0_m3_M1_X0_Y0_1 net_m0_m3_M1_X0_Y0_diff net_m0_m3_M1_X0_Y0_G net_m0_m3_M1_X0_Y0_S gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m0_m3_M2_X1_Y0_0 net_m0_m3_M2_X1_Y0_D net_m0_m3_M2_X1_Y0_G net_m0_m3_M2_X1_Y0_diff gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12
x_m0_m3_M2_X1_Y0_1 net_m0_m3_M2_X1_Y0_diff net_m0_m3_M2_X1_Y0_G net_m0_m3_M2_X1_Y0_S gnd! nmos_rvt w=2.7e-07 l=2e-08 nfin=12

**connections
v_vdd_inject vdd! vdd_M4_3040_336 0
v_id_inject id id_M3_640_252 0
v_vinp_inject vinp vinp_M5_1440_0 0
v_vinn_inject vinn vinn_M2_2400_504 0
v_vout_probe vout_M4_2440_252 vout 0
v_vss_inject 0 vss_M3_560_132 0
v_net10_probe net10 net10_M4_960_168 0
v_net8_probe net8 net8_M4_3680_420 0

**testbench
v2 vinp 0 DC 675e-3 AC 0.5 180 SIN(675e-3 .002 1k 0 0 180)
v1 vinn 0 DC 675e-3 AC 0.5     SIN(675e-3 .002 1k 0 0   0)
v0 vdd! 0 1.0
i5 vdd! id 40e-6
cload vout 0 350e-15

*.OP

*.PRINT DC v(vout) v(id) v(vinp) v(vinn) id(x_m5_m4_M2_X1_Y0_0:mn) id(x_m5_m4_M2_X1_Y0_1:mn) id(x_m5_m4_M1_X0_Y0_0:mn) id(x_m5_m4_M1_X0_Y0_1:mn)

.AC DEC 100 1.0 1e11

.PRINT AC vdb(vout) vm(vout)

*.tran 10n 5m
*.PRINT TRAN v(vout) v(vinp) v(vinn) v(id) v(net10) v(net8) id(x_m5_m4_M2_X1_Y0_0:mn)
*.OPTIONS OUTPUT INITIAL_INTERVAL=1u
*.OPTIONS TIMEINT RELTOL=1e-4 ABSTOL=1e-8

*.MEASURE TRAN vout_max MAX v(vout)
*.MEASURE TRAN vout_min MIN v(vout)
*.MEASURE TRAN vout_pp  PP  v(vout)

.END

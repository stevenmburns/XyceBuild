
*
* Short channel models from CMOS Circuit Design, Layout, and Simulation,
* 50nm BSIM4 models VDD=1V, see CMOSedu.com
*
.model  N_50n  nmos  level = 54
+binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 0          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0          
+tnom    = 27           toxe    = 1.4e-009     toxp    = 7e-010       toxm    = 1.4e-009   
+epsrox  = 3.9          wint    = 5e-009       lint    = 1.2e-008   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 1.4e-009   
+vth0    = 0.22         k1      = 0.35         k2      = 0.05         k3      = 0          
+k3b     = 0            w0      = 2.5e-006     dvt0    = 2.8          dvt1    = 0.52       
+dvt2    = -0.032       dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 2            minv    = 0.05         voffl   = 0            dvtp0   = 1e-007     
+dvtp1   = 0.05         lpe0    = 5.75e-008    lpeb    = 2.3e-010     xj      = 2e-008     
+ngate   = 5e+020       ndep    = 2.8e+018     nsd     = 1e+020       phin    = 0          
+cdsc    = 0.0002       cdscb   = 0            cdscd   = 0            cit     = 0          
+voff    = -0.15        nfactor = 1.2          eta0    = 0.15         etab    = 0          
+vfb     = -0.55        u0      = 0.032        ua      = 1.6e-010     ub      = 1.1e-017   
+uc      = -3e-011      vsat    = 1.1e+005     a0      = 2            ags     = 1e-020     
+a1      = 0            a2      = 1            b0      = -1e-020      b1      = 0          
+keta    = 0.04         dwg     = 0            dwb     = 0            pclm    = 0.18       
+pdiblc1 = 0.028        pdiblc2 = 0.022        pdiblcb = -0.005       drout   = 0.45       
+pvag    = 1e-020       delta   = 0.01         pscbe1  = 8.14e+008    pscbe2  = 1e-007     
+fprout  = 0.2          pdits   = 0.2          pditsd  = 0.23         pditsl  = 2.3e+006   
+rsh     = 3            rdsw    = 150          rsw     = 150          rdw     = 150        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 0          
+prwb    = 6.8e-011     wr      = 1            alpha0  = 0.074        alpha1  = 0.005      
+beta0   = 30           agidl   = 0.0002       bgidl   = 2.1e+009     cgidl   = 0.0002     
+egidl   = 0.8          
+aigbacc = 0.012        bigbacc = 0.0028       cigbacc = 0.002
+nigbacc = 1            aigbinv = 0.014        bigbinv = 0.004        cigbinv = 0.004
+eigbinv = 1.1          nigbinv = 3            aigc    = 0.017        bigc    = 0.0028
+cigc    = 0.002        aigsd   = 0.017        bigsd   = 0.0028       cigsd   = 0.002
+nigc    = 1            poxedge = 1            pigcd   = 1            ntox    = 1
+xrcrg1  = 12           xrcrg2  = 5          
+cgso    = 6.238e-010   cgdo    = 6.238e-010   cgbo    = 2.56e-011    cgdl    = 2.495e-10     
+cgsl    = 2.495e-10    ckappas = 0.02         ckappad = 0.02         acde    = 1          
+moin    = 15           noff    = 0.9          voffcv  = 0.02       
+kt1     = -0.21        kt1l    = 0.0           kt2     = -0.042        ute     = -1.5
+ua1     = 1e-009       ub1     = -3.5e-019     uc1     = 0             prt     = 0
+at      = 53000
+fnoimod = 1            tnoimod = 0          
+jss     = 0.0001       jsws    = 1e-011       jswgs   = 1e-010       njs     = 1          
+ijthsfwd= 0.01         ijthsrev= 0.001        bvs     = 10           xjbvs   = 1          
+jsd     = 0.0001       jswd    = 1e-011       jswgd   = 1e-010       njd     = 1          
+ijthdfwd= 0.01         ijthdrev= 0.001        bvd     = 10           xjbvd   = 1          
+pbs     = 1            cjs     = 0.0005       mjs     = 0.5          pbsws   = 1          
+cjsws   = 5e-010       mjsws   = 0.33         pbswgs  = 1            cjswgs  = 5e-010     
+mjswgs  = 0.33         pbd     = 1            cjd     = 0.0005       mjd     = 0.5        
+pbswd   = 1            cjswd   = 5e-010       mjswd   = 0.33         pbswgd  = 1          
+cjswgd  = 5e-010       mjswgd  = 0.33         tpb     = 0.005        tcj     = 0.001      
+tpbsw   = 0.005        tcjsw   = 0.001        tpbswg  = 0.005        tcjswg  = 0.001      
+xtis    = 3            xtid    = 3          
+dmcg    = 0e-006       dmci    = 0e-006       dmdg    = 0e-006       dmcgt   = 0e-007     
+dwj     = 0e-008     	xgw     = 0e-007       xgl     = 0e-008     
+rshg    = 0.4          gbmin   = 1e-010       rbpb    = 5            rbpd    = 15         
+rbps    = 15           rbdb    = 15           rbsb    = 15           ngcon   = 1
*
.model  P_50n  pmos  level = 54
+binunit = 1            paramchk= 1            mobmod  = 0          
+capmod  = 2            igcmod  = 1            igbmod  = 1            geomod  = 0          
+diomod  = 1            rdsmod  = 0            rbodymod= 1            rgatemod= 1          
+permod  = 1            acnqsmod= 0            trnqsmod= 0          
+tnom    = 27           toxe    = 1.4e-009     toxp    = 7e-010       toxm    = 1.4e-009   
+epsrox  = 3.9          wint    = 5e-009       lint    = 1.2e-008   
+ll      = 0            wl      = 0            lln     = 1            wln     = 1          
+lw      = 0            ww      = 0            lwn     = 1            wwn     = 1          
+lwl     = 0            wwl     = 0            xpart   = 0            toxref  = 1.4e-009   
+vth0    = -0.22        k1      = 0.39         k2      = 0.05         k3      = 0          
+k3b     = 0            w0      = 2.5e-006     dvt0    = 3.9          dvt1    = 0.635        
+dvt2    = -0.032       dvt0w   = 0            dvt1w   = 0            dvt2w   = 0          
+dsub    = 0.7          minv    = 0.05         voffl   = 0            dvtp0   = 0.5e-008     
+dvtp1   = 0.05         lpe0    = 5.75e-008    lpeb    = 2.3e-010     xj      = 2e-008     
+ngate   = 5e+020       ndep    = 2.8e+018     nsd     = 1e+020       phin    = 0          
+cdsc    = 0.000258     cdscb   = 0            cdscd   = 6.1e-008     cit     = 0          
+voff    = -0.15        nfactor = 2            eta0    = 0.15         etab    = 0          
+vfb     = 0.55         u0      = 0.0095       ua      = 1.6e-009     ub      = 8e-018     
+uc      = 4.6e-013     vsat    = 90000        a0      = 1.2          ags     = 1e-020     
+a1      = 0            a2      = 1            b0      = -1e-020      b1      = 0          
+keta    = -0.047       dwg     = 0            dwb     = 0            pclm    = 0.55       
+pdiblc1 = 0.03         pdiblc2 = 0.0055       pdiblcb = 3.4e-008     drout   = 0.56       
+pvag    = 1e-020       delta   = 0.014        pscbe1  = 8.14e+008    pscbe2  = 9.58e-007  
+fprout  = 0.2          pdits   = 0.2          pditsd  = 0.23         pditsl  = 2.3e+006   
+rsh     = 3            rdsw    = 250          rsw     = 160          rdw     = 160        
+rdswmin = 0            rdwmin  = 0            rswmin  = 0            prwg    = 3.22e-008  
+prwb    = 6.8e-011     wr      = 1            alpha0  = 0.074        alpha1  = 0.005      
+beta0   = 30           agidl   = 0.0002       bgidl   = 2.1e+009     cgidl   = 0.0002     
+egidl   = 0.8          
+aigbacc = 0.012        bigbacc = 0.0028       cigbacc = 0.002
+nigbacc = 1            aigbinv = 0.014        bigbinv = 0.004        cigbinv = 0.004
+eigbinv = 1.1          nigbinv = 3            aigc    = 0.69         bigc    = 0.0012
+cigc    = 0.0008       aigsd   = 0.0087       bigsd   = 0.0012       cigsd   = 0.0008
+nigc    = 1            poxedge = 1            pigcd   = 1            ntox    = 1
+xrcrg1  = 12           xrcrg2  = 5          
+cgso    = 7.43e-010    cgdo    = 7.43e-010    cgbo    = 2.56e-011    cgdl    = 1e-014     
+cgsl    = 1e-014       ckappas = 0.5          ckappad = 0.5          acde    = 1          
+moin    = 15           noff    = 0.9          voffcv  = 0.02       
+kt1     = -0.19        kt1l    = 0            kt2     = -0.052        ute     = -1.5
+ua1     = -1e-009      ub1     = 2e-018       uc1     = 0             prt     = 0
+at      = 33000
+fnoimod = 1            tnoimod = 0          
+jss     = 0.0001       jsws    = 1e-011       jswgs   = 1e-010       njs     = 1          
+ijthsfwd= 0.01         ijthsrev= 0.001        bvs     = 10           xjbvs   = 1          
+jsd     = 0.0001       jswd    = 1e-011       jswgd   = 1e-010       njd     = 1          
+ijthdfwd= 0.01         ijthdrev= 0.001        bvd     = 10           xjbvd   = 1          
+pbs     = 1            cjs     = 0.0005       mjs     = 0.5          pbsws   = 1          
+cjsws   = 5e-010       mjsws   = 0.33         pbswgs  = 1            cjswgs  = 5e-010     
+mjswgs  = 0.33         pbd     = 1            cjd     = 0.0005       mjd     = 0.5        
+pbswd   = 1            cjswd   = 5e-010       mjswd   = 0.33         pbswgd  = 1          
+cjswgd  = 5e-010       mjswgd  = 0.33         tpb     = 0.005        tcj     = 0.001      
+tpbsw   = 0.005        tcjsw   = 0.001        tpbswg  = 0.005        tcjswg  = 0.001      
+xtis    = 3            xtid    = 3          
+dmcg    = 0e-006       dmci    = 0e-006       dmdg    = 0e-006       dmcgt   = 0e-007     
+dwj     = 0e-008     	xgw     = 0e-007       xgl     = 0e-008     
+rshg    = 0.4          gbmin   = 1e-010       rbpb    = 5            rbpd    = 15         
+rbps    = 15           rbdb    = 15           rbsb    = 15           ngcon   = 1   


.MODEL NMOS NMOS
.MODEL PMOS PMOS

.GLOBAL vdd!

*.TEMP 25.0

*.OPTION INGOLD=2 ARTIST=2 PSF=2 MEASOUT=1 PARHIER=LOCAL PROBE=0 MARCH=2 ACCURACY=1 POST

.SUBCKT NMOS d g s b PARAMS: w=270e-9 l=20e-9 nfin=10
.param width={nfin*100n}
.param length={50n}
.param perimeter={3*length}
.param area={1.5*length*width}

mn d g s b N_50n L={length} W={width} PD={perimeter} AD={area}
.ENDS

.SUBCKT PMOS d g s b PARAMS: w=270e-9 l=20e-9 nfin=10
.param width={nfin*100n}
.param length={2*50n}
.param perimeter={3*length}
.param area={1.5*length*width}

mp d g s b P_50n L={length} W={width} PD={perimeter} AD={area}
.ENDS

r0 net8_M1_3840_132 net8_M1_3840_212 8.0
c0 net8_M1_3840_132 0 0.008f
c1 net8_M1_3840_212 0 0.008f
r1 net8_M1_3840_212 net8_M1_3840_252 4.0
c2 net8_M1_3840_212 0 0.004f
c3 net8_M1_3840_252 0 0.004f
r2 net8_M1_3840_252 net8_M1_3840_332 8.0
c4 net8_M1_3840_252 0 0.008f
c5 net8_M1_3840_332 0 0.008f
r3 net8_M1_3840_332 net8_M1_3840_412 8.0
c6 net8_M1_3840_332 0 0.008f
c7 net8_M1_3840_412 0 0.008f
r4 net8_M1_3840_412 net8_M1_3840_420 0.8
c8 net8_M1_3840_412 0 0.0008f
c9 net8_M1_3840_420 0 0.0008f
r5 net8_M1_3840_168 net8_M1_3840_248 8.0
c10 net8_M1_3840_168 0 0.008f
c11 net8_M1_3840_248 0 0.008f
r6 net8_M1_3840_248 net8_M1_3840_328 8.0
c12 net8_M1_3840_248 0 0.008f
c13 net8_M1_3840_328 0 0.008f
r7 net8_M1_3840_328 net8_M1_3840_408 8.0
c14 net8_M1_3840_328 0 0.008f
c15 net8_M1_3840_408 0 0.008f
r8 net8_M1_3840_408 net8_M1_3840_488 8.0
c16 net8_M1_3840_408 0 0.008f
c17 net8_M1_3840_488 0 0.008f
r9 net8_M1_3840_488 net8_M1_3840_568 8.0
c18 net8_M1_3840_488 0 0.008f
c19 net8_M1_3840_568 0 0.008f
r10 net8_M1_3840_568 net8_M1_3840_648 8.0
c20 net8_M1_3840_568 0 0.008f
c21 net8_M1_3840_648 0 0.008f
r11 net8_M1_3840_648 net8_M1_3840_728 8.0
c22 net8_M1_3840_648 0 0.008f
c23 net8_M1_3840_728 0 0.008f
r12 net8_M1_3840_728 net8_M1_3840_792 6.4
c24 net8_M1_3840_728 0 0.0064f
c25 net8_M1_3840_792 0 0.0064f
r13 vdd_M1_3920_132 vdd_M1_3920_168 3.5999999999999996
c26 vdd_M1_3920_132 0 0.0036f
c27 vdd_M1_3920_168 0 0.0036f
r14 vdd_M1_3920_168 vdd_M1_3920_248 8.0
c28 vdd_M1_3920_168 0 0.008f
c29 vdd_M1_3920_248 0 0.008f
r15 vdd_M1_3920_248 vdd_M1_3920_328 8.0
c30 vdd_M1_3920_248 0 0.008f
c31 vdd_M1_3920_328 0 0.008f
r16 vdd_M1_3920_328 vdd_M1_3920_336 0.8
c32 vdd_M1_3920_328 0 0.0008f
c33 vdd_M1_3920_336 0 0.0008f
r17 vdd_M1_3920_336 vdd_M1_3920_416 8.0
c34 vdd_M1_3920_336 0 0.008f
c35 vdd_M1_3920_416 0 0.008f
r18 vdd_M1_3920_416 vdd_M1_3920_462 4.6
c36 vdd_M1_3920_416 0 0.0046f
c37 vdd_M1_3920_462 0 0.0046f
r19 vdd_M1_3920_462 vdd_M1_3920_542 8.0
c38 vdd_M1_3920_462 0 0.008f
c39 vdd_M1_3920_542 0 0.008f
r20 vdd_M1_3920_542 vdd_M1_3920_588 4.6
c40 vdd_M1_3920_542 0 0.0046f
c41 vdd_M1_3920_588 0 0.0046f
r21 vdd_M1_3920_588 vdd_M1_3920_668 8.0
c42 vdd_M1_3920_588 0 0.008f
c43 vdd_M1_3920_668 0 0.008f
r22 vdd_M1_3920_668 vdd_M1_3920_748 8.0
c44 vdd_M1_3920_668 0 0.008f
c45 vdd_M1_3920_748 0 0.008f
r23 vdd_M1_3920_748 vdd_M1_3920_792 4.3999999999999995
c46 vdd_M1_3920_748 0 0.0044f
c47 vdd_M1_3920_792 0 0.0044f
r24 net8_M1_3760_132 net8_M1_3760_212 8.0
c48 net8_M1_3760_132 0 0.008f
c49 net8_M1_3760_212 0 0.008f
r25 net8_M1_3760_212 net8_M1_3760_252 4.0
c50 net8_M1_3760_212 0 0.004f
c51 net8_M1_3760_252 0 0.004f
r26 net8_M1_3760_252 net8_M1_3760_332 8.0
c52 net8_M1_3760_252 0 0.008f
c53 net8_M1_3760_332 0 0.008f
r27 net8_M1_3760_332 net8_M1_3760_412 8.0
c54 net8_M1_3760_332 0 0.008f
c55 net8_M1_3760_412 0 0.008f
r28 net8_M1_3760_412 net8_M1_3760_420 0.8
c56 net8_M1_3760_412 0 0.0008f
c57 net8_M1_3760_420 0 0.0008f
r29 net8_M1_3760_336 net8_M1_3760_416 8.0
c58 net8_M1_3760_336 0 0.008f
c59 net8_M1_3760_416 0 0.008f
r30 net8_M1_3760_416 net8_M1_3760_462 4.6
c60 net8_M1_3760_416 0 0.0046f
c61 net8_M1_3760_462 0 0.0046f
r31 net8_M1_3760_462 net8_M1_3760_542 8.0
c62 net8_M1_3760_462 0 0.008f
c63 net8_M1_3760_542 0 0.008f
r32 net8_M1_3760_542 net8_M1_3760_588 4.6
c64 net8_M1_3760_542 0 0.0046f
c65 net8_M1_3760_588 0 0.0046f
r33 net8_M1_3760_588 net8_M1_3760_668 8.0
c66 net8_M1_3760_588 0 0.008f
c67 net8_M1_3760_668 0 0.008f
r34 net8_M1_3760_668 net8_M1_3760_748 8.0
c68 net8_M1_3760_668 0 0.008f
c69 net8_M1_3760_748 0 0.008f
r35 net8_M1_3760_748 net8_M1_3760_792 4.3999999999999995
c70 net8_M1_3760_748 0 0.0044f
c71 net8_M1_3760_792 0 0.0044f
r36 net8_M1_3120_132 net8_M1_3120_212 8.0
c72 net8_M1_3120_132 0 0.008f
c73 net8_M1_3120_212 0 0.008f
r37 net8_M1_3120_212 net8_M1_3120_292 8.0
c74 net8_M1_3120_212 0 0.008f
c75 net8_M1_3120_292 0 0.008f
r38 net8_M1_3120_292 net8_M1_3120_336 4.3999999999999995
c76 net8_M1_3120_292 0 0.0044f
c77 net8_M1_3120_336 0 0.0044f
r39 net8_M1_3120_336 net8_M1_3120_416 8.0
c78 net8_M1_3120_336 0 0.008f
c79 net8_M1_3120_416 0 0.008f
r40 net8_M1_3120_416 net8_M1_3120_496 8.0
c80 net8_M1_3120_416 0 0.008f
c81 net8_M1_3120_496 0 0.008f
r41 net8_M1_3120_496 net8_M1_3120_576 8.0
c82 net8_M1_3120_496 0 0.008f
c83 net8_M1_3120_576 0 0.008f
r42 net8_M1_3120_576 net8_M1_3120_588 1.2
c84 net8_M1_3120_576 0 0.0012000000000000001f
c85 net8_M1_3120_588 0 0.0012000000000000001f
r43 net8_M1_3120_168 net8_M1_3120_248 8.0
c86 net8_M1_3120_168 0 0.008f
c87 net8_M1_3120_248 0 0.008f
r44 net8_M1_3120_248 net8_M1_3120_328 8.0
c88 net8_M1_3120_248 0 0.008f
c89 net8_M1_3120_328 0 0.008f
r45 net8_M1_3120_328 net8_M1_3120_408 8.0
c90 net8_M1_3120_328 0 0.008f
c91 net8_M1_3120_408 0 0.008f
r46 net8_M1_3120_408 net8_M1_3120_488 8.0
c92 net8_M1_3120_408 0 0.008f
c93 net8_M1_3120_488 0 0.008f
r47 net8_M1_3120_488 net8_M1_3120_568 8.0
c94 net8_M1_3120_488 0 0.008f
c95 net8_M1_3120_568 0 0.008f
r48 net8_M1_3120_568 net8_M1_3120_648 8.0
c96 net8_M1_3120_568 0 0.008f
c97 net8_M1_3120_648 0 0.008f
r49 net8_M1_3120_648 net8_M1_3120_728 8.0
c98 net8_M1_3120_648 0 0.008f
c99 net8_M1_3120_728 0 0.008f
r50 net8_M1_3120_728 net8_M1_3120_792 6.4
c100 net8_M1_3120_728 0 0.0064f
c101 net8_M1_3120_792 0 0.0064f
r51 vdd_M1_3200_132 vdd_M1_3200_168 3.5999999999999996
c102 vdd_M1_3200_132 0 0.0036f
c103 vdd_M1_3200_168 0 0.0036f
r52 vdd_M1_3200_168 vdd_M1_3200_248 8.0
c104 vdd_M1_3200_168 0 0.008f
c105 vdd_M1_3200_248 0 0.008f
r53 vdd_M1_3200_248 vdd_M1_3200_328 8.0
c106 vdd_M1_3200_248 0 0.008f
c107 vdd_M1_3200_328 0 0.008f
r54 vdd_M1_3200_328 vdd_M1_3200_408 8.0
c108 vdd_M1_3200_328 0 0.008f
c109 vdd_M1_3200_408 0 0.008f
r55 vdd_M1_3200_408 vdd_M1_3200_420 1.2
c110 vdd_M1_3200_408 0 0.0012000000000000001f
c111 vdd_M1_3200_420 0 0.0012000000000000001f
r56 vdd_M1_3200_336 vdd_M1_3200_416 8.0
c112 vdd_M1_3200_336 0 0.008f
c113 vdd_M1_3200_416 0 0.008f
r57 vdd_M1_3200_416 vdd_M1_3200_462 4.6
c114 vdd_M1_3200_416 0 0.0046f
c115 vdd_M1_3200_462 0 0.0046f
r58 vdd_M1_3200_462 vdd_M1_3200_542 8.0
c116 vdd_M1_3200_462 0 0.008f
c117 vdd_M1_3200_542 0 0.008f
r59 vdd_M1_3200_542 vdd_M1_3200_588 4.6
c118 vdd_M1_3200_542 0 0.0046f
c119 vdd_M1_3200_588 0 0.0046f
r60 vdd_M1_3200_588 vdd_M1_3200_668 8.0
c120 vdd_M1_3200_588 0 0.008f
c121 vdd_M1_3200_668 0 0.008f
r61 vdd_M1_3200_668 vdd_M1_3200_748 8.0
c122 vdd_M1_3200_668 0 0.008f
c123 vdd_M1_3200_748 0 0.008f
r62 vdd_M1_3200_748 vdd_M1_3200_792 4.3999999999999995
c124 vdd_M1_3200_748 0 0.0044f
c125 vdd_M1_3200_792 0 0.0044f
r63 vout_M1_3040_132 vout_M1_3040_212 8.0
c126 vout_M1_3040_132 0 0.008f
c127 vout_M1_3040_212 0 0.008f
r64 vout_M1_3040_212 vout_M1_3040_252 4.0
c128 vout_M1_3040_212 0 0.004f
c129 vout_M1_3040_252 0 0.004f
r65 vout_M1_3040_252 vout_M1_3040_332 8.0
c130 vout_M1_3040_252 0 0.008f
c131 vout_M1_3040_332 0 0.008f
r66 vout_M1_3040_332 vout_M1_3040_412 8.0
c132 vout_M1_3040_332 0 0.008f
c133 vout_M1_3040_412 0 0.008f
r67 vout_M1_3040_412 vout_M1_3040_492 8.0
c134 vout_M1_3040_412 0 0.008f
c135 vout_M1_3040_492 0 0.008f
r68 vout_M1_3040_492 vout_M1_3040_504 1.2
c136 vout_M1_3040_492 0 0.0012000000000000001f
c137 vout_M1_3040_504 0 0.0012000000000000001f
r69 vout_M1_3040_336 vout_M1_3040_416 8.0
c138 vout_M1_3040_336 0 0.008f
c139 vout_M1_3040_416 0 0.008f
r70 vout_M1_3040_416 vout_M1_3040_462 4.6
c140 vout_M1_3040_416 0 0.0046f
c141 vout_M1_3040_462 0 0.0046f
r71 vout_M1_3040_462 vout_M1_3040_542 8.0
c142 vout_M1_3040_462 0 0.008f
c143 vout_M1_3040_542 0 0.008f
r72 vout_M1_3040_542 vout_M1_3040_588 4.6
c144 vout_M1_3040_542 0 0.0046f
c145 vout_M1_3040_588 0 0.0046f
r73 vout_M1_3040_588 vout_M1_3040_668 8.0
c146 vout_M1_3040_588 0 0.008f
c147 vout_M1_3040_668 0 0.008f
r74 vout_M1_3040_668 vout_M1_3040_748 8.0
c148 vout_M1_3040_668 0 0.008f
c149 vout_M1_3040_748 0 0.008f
r75 vout_M1_3040_748 vout_M1_3040_792 4.3999999999999995
c150 vout_M1_3040_748 0 0.0044f
c151 vout_M1_3040_792 0 0.0044f
r76 id_M1_400_132 id_M1_400_212 8.0
c152 id_M1_400_132 0 0.008f
c153 id_M1_400_212 0 0.008f
r77 id_M1_400_212 id_M1_400_252 4.0
c154 id_M1_400_212 0 0.004f
c155 id_M1_400_252 0 0.004f
r78 id_M1_400_252 id_M1_400_332 8.0
c156 id_M1_400_252 0 0.008f
c157 id_M1_400_332 0 0.008f
r79 id_M1_400_332 id_M1_400_412 8.0
c158 id_M1_400_332 0 0.008f
c159 id_M1_400_412 0 0.008f
r80 id_M1_400_412 id_M1_400_492 8.0
c160 id_M1_400_412 0 0.008f
c161 id_M1_400_492 0 0.008f
r81 id_M1_400_492 id_M1_400_504 1.2
c162 id_M1_400_492 0 0.0012000000000000001f
c163 id_M1_400_504 0 0.0012000000000000001f
r82 id_M1_400_168 id_M1_400_248 8.0
c164 id_M1_400_168 0 0.008f
c165 id_M1_400_248 0 0.008f
r83 id_M1_400_248 id_M1_400_328 8.0
c166 id_M1_400_248 0 0.008f
c167 id_M1_400_328 0 0.008f
r84 id_M1_400_328 id_M1_400_408 8.0
c168 id_M1_400_328 0 0.008f
c169 id_M1_400_408 0 0.008f
r85 id_M1_400_408 id_M1_400_488 8.0
c170 id_M1_400_408 0 0.008f
c171 id_M1_400_488 0 0.008f
r86 id_M1_400_488 id_M1_400_568 8.0
c172 id_M1_400_488 0 0.008f
c173 id_M1_400_568 0 0.008f
r87 id_M1_400_568 id_M1_400_648 8.0
c174 id_M1_400_568 0 0.008f
c175 id_M1_400_648 0 0.008f
r88 id_M1_400_648 id_M1_400_728 8.0
c176 id_M1_400_648 0 0.008f
c177 id_M1_400_728 0 0.008f
r89 id_M1_400_728 id_M1_400_792 6.4
c178 id_M1_400_728 0 0.0064f
c179 id_M1_400_792 0 0.0064f
r90 vss_M1_320_132 vss_M1_320_168 3.5999999999999996
c180 vss_M1_320_132 0 0.0036f
c181 vss_M1_320_168 0 0.0036f
r91 vss_M1_320_168 vss_M1_320_248 8.0
c182 vss_M1_320_168 0 0.008f
c183 vss_M1_320_248 0 0.008f
r92 vss_M1_320_248 vss_M1_320_328 8.0
c184 vss_M1_320_248 0 0.008f
c185 vss_M1_320_328 0 0.008f
r93 vss_M1_320_328 vss_M1_320_408 8.0
c186 vss_M1_320_328 0 0.008f
c187 vss_M1_320_408 0 0.008f
r94 vss_M1_320_408 vss_M1_320_420 1.2
c188 vss_M1_320_408 0 0.0012000000000000001f
c189 vss_M1_320_420 0 0.0012000000000000001f
r95 vss_M1_320_336 vss_M1_320_416 8.0
c190 vss_M1_320_336 0 0.008f
c191 vss_M1_320_416 0 0.008f
r96 vss_M1_320_416 vss_M1_320_462 4.6
c192 vss_M1_320_416 0 0.0046f
c193 vss_M1_320_462 0 0.0046f
r97 vss_M1_320_462 vss_M1_320_542 8.0
c194 vss_M1_320_462 0 0.008f
c195 vss_M1_320_542 0 0.008f
r98 vss_M1_320_542 vss_M1_320_588 4.6
c196 vss_M1_320_542 0 0.0046f
c197 vss_M1_320_588 0 0.0046f
r99 vss_M1_320_588 vss_M1_320_668 8.0
c198 vss_M1_320_588 0 0.008f
c199 vss_M1_320_668 0 0.008f
r100 vss_M1_320_668 vss_M1_320_748 8.0
c200 vss_M1_320_668 0 0.008f
c201 vss_M1_320_748 0 0.008f
r101 vss_M1_320_748 vss_M1_320_792 4.3999999999999995
c202 vss_M1_320_748 0 0.0044f
c203 vss_M1_320_792 0 0.0044f
r102 id_M1_480_132 id_M1_480_212 8.0
c204 id_M1_480_132 0 0.008f
c205 id_M1_480_212 0 0.008f
r103 id_M1_480_212 id_M1_480_252 4.0
c206 id_M1_480_212 0 0.004f
c207 id_M1_480_252 0 0.004f
r104 id_M1_480_252 id_M1_480_332 8.0
c208 id_M1_480_252 0 0.008f
c209 id_M1_480_332 0 0.008f
r105 id_M1_480_332 id_M1_480_412 8.0
c210 id_M1_480_332 0 0.008f
c211 id_M1_480_412 0 0.008f
r106 id_M1_480_412 id_M1_480_492 8.0
c212 id_M1_480_412 0 0.008f
c213 id_M1_480_492 0 0.008f
r107 id_M1_480_492 id_M1_480_504 1.2
c214 id_M1_480_492 0 0.0012000000000000001f
c215 id_M1_480_504 0 0.0012000000000000001f
r108 id_M1_480_336 id_M1_480_416 8.0
c216 id_M1_480_336 0 0.008f
c217 id_M1_480_416 0 0.008f
r109 id_M1_480_416 id_M1_480_462 4.6
c218 id_M1_480_416 0 0.0046f
c219 id_M1_480_462 0 0.0046f
r110 id_M1_480_462 id_M1_480_542 8.0
c220 id_M1_480_462 0 0.008f
c221 id_M1_480_542 0 0.008f
r111 id_M1_480_542 id_M1_480_588 4.6
c222 id_M1_480_542 0 0.0046f
c223 id_M1_480_588 0 0.0046f
r112 id_M1_480_588 id_M1_480_668 8.0
c224 id_M1_480_588 0 0.008f
c225 id_M1_480_668 0 0.008f
r113 id_M1_480_668 id_M1_480_748 8.0
c226 id_M1_480_668 0 0.008f
c227 id_M1_480_748 0 0.008f
r114 id_M1_480_748 id_M1_480_792 4.3999999999999995
c228 id_M1_480_748 0 0.0044f
c229 id_M1_480_792 0 0.0044f
r115 id_M1_1040_132 id_M1_1040_212 8.0
c230 id_M1_1040_132 0 0.008f
c231 id_M1_1040_212 0 0.008f
r116 id_M1_1040_212 id_M1_1040_252 4.0
c232 id_M1_1040_212 0 0.004f
c233 id_M1_1040_252 0 0.004f
r117 id_M1_1040_252 id_M1_1040_332 8.0
c234 id_M1_1040_252 0 0.008f
c235 id_M1_1040_332 0 0.008f
r118 id_M1_1040_332 id_M1_1040_412 8.0
c236 id_M1_1040_332 0 0.008f
c237 id_M1_1040_412 0 0.008f
r119 id_M1_1040_412 id_M1_1040_492 8.0
c238 id_M1_1040_412 0 0.008f
c239 id_M1_1040_492 0 0.008f
r120 id_M1_1040_492 id_M1_1040_504 1.2
c240 id_M1_1040_492 0 0.0012000000000000001f
c241 id_M1_1040_504 0 0.0012000000000000001f
r121 id_M1_1040_168 id_M1_1040_248 8.0
c242 id_M1_1040_168 0 0.008f
c243 id_M1_1040_248 0 0.008f
r122 id_M1_1040_248 id_M1_1040_328 8.0
c244 id_M1_1040_248 0 0.008f
c245 id_M1_1040_328 0 0.008f
r123 id_M1_1040_328 id_M1_1040_408 8.0
c246 id_M1_1040_328 0 0.008f
c247 id_M1_1040_408 0 0.008f
r124 id_M1_1040_408 id_M1_1040_488 8.0
c248 id_M1_1040_408 0 0.008f
c249 id_M1_1040_488 0 0.008f
r125 id_M1_1040_488 id_M1_1040_568 8.0
c250 id_M1_1040_488 0 0.008f
c251 id_M1_1040_568 0 0.008f
r126 id_M1_1040_568 id_M1_1040_648 8.0
c252 id_M1_1040_568 0 0.008f
c253 id_M1_1040_648 0 0.008f
r127 id_M1_1040_648 id_M1_1040_728 8.0
c254 id_M1_1040_648 0 0.008f
c255 id_M1_1040_728 0 0.008f
r128 id_M1_1040_728 id_M1_1040_792 6.4
c256 id_M1_1040_728 0 0.0064f
c257 id_M1_1040_792 0 0.0064f
r129 vss_M1_960_132 vss_M1_960_168 3.5999999999999996
c258 vss_M1_960_132 0 0.0036f
c259 vss_M1_960_168 0 0.0036f
r130 vss_M1_960_168 vss_M1_960_248 8.0
c260 vss_M1_960_168 0 0.008f
c261 vss_M1_960_248 0 0.008f
r131 vss_M1_960_248 vss_M1_960_328 8.0
c262 vss_M1_960_248 0 0.008f
c263 vss_M1_960_328 0 0.008f
r132 vss_M1_960_328 vss_M1_960_408 8.0
c264 vss_M1_960_328 0 0.008f
c265 vss_M1_960_408 0 0.008f
r133 vss_M1_960_408 vss_M1_960_420 1.2
c266 vss_M1_960_408 0 0.0012000000000000001f
c267 vss_M1_960_420 0 0.0012000000000000001f
r134 vss_M1_960_336 vss_M1_960_416 8.0
c268 vss_M1_960_336 0 0.008f
c269 vss_M1_960_416 0 0.008f
r135 vss_M1_960_416 vss_M1_960_462 4.6
c270 vss_M1_960_416 0 0.0046f
c271 vss_M1_960_462 0 0.0046f
r136 vss_M1_960_462 vss_M1_960_542 8.0
c272 vss_M1_960_462 0 0.008f
c273 vss_M1_960_542 0 0.008f
r137 vss_M1_960_542 vss_M1_960_588 4.6
c274 vss_M1_960_542 0 0.0046f
c275 vss_M1_960_588 0 0.0046f
r138 vss_M1_960_588 vss_M1_960_668 8.0
c276 vss_M1_960_588 0 0.008f
c277 vss_M1_960_668 0 0.008f
r139 vss_M1_960_668 vss_M1_960_748 8.0
c278 vss_M1_960_668 0 0.008f
c279 vss_M1_960_748 0 0.008f
r140 vss_M1_960_748 vss_M1_960_792 4.3999999999999995
c280 vss_M1_960_748 0 0.0044f
c281 vss_M1_960_792 0 0.0044f
r141 net10_M1_1120_132 net10_M1_1120_212 8.0
c282 net10_M1_1120_132 0 0.008f
c283 net10_M1_1120_212 0 0.008f
r142 net10_M1_1120_212 net10_M1_1120_292 8.0
c284 net10_M1_1120_212 0 0.008f
c285 net10_M1_1120_292 0 0.008f
r143 net10_M1_1120_292 net10_M1_1120_336 4.3999999999999995
c286 net10_M1_1120_292 0 0.0044f
c287 net10_M1_1120_336 0 0.0044f
r144 net10_M1_1120_336 net10_M1_1120_416 8.0
c288 net10_M1_1120_336 0 0.008f
c289 net10_M1_1120_416 0 0.008f
r145 net10_M1_1120_416 net10_M1_1120_496 8.0
c290 net10_M1_1120_416 0 0.008f
c291 net10_M1_1120_496 0 0.008f
r146 net10_M1_1120_496 net10_M1_1120_576 8.0
c292 net10_M1_1120_496 0 0.008f
c293 net10_M1_1120_576 0 0.008f
r147 net10_M1_1120_576 net10_M1_1120_588 1.2
c294 net10_M1_1120_576 0 0.0012000000000000001f
c295 net10_M1_1120_588 0 0.0012000000000000001f
r148 net10_M1_1120_462 net10_M1_1120_542 8.0
c296 net10_M1_1120_462 0 0.008f
c297 net10_M1_1120_542 0 0.008f
r149 net10_M1_1120_542 net10_M1_1120_622 8.0
c298 net10_M1_1120_542 0 0.008f
c299 net10_M1_1120_622 0 0.008f
r150 net10_M1_1120_622 net10_M1_1120_702 8.0
c300 net10_M1_1120_622 0 0.008f
c301 net10_M1_1120_702 0 0.008f
r151 net10_M1_1120_702 net10_M1_1120_782 8.0
c302 net10_M1_1120_702 0 0.008f
c303 net10_M1_1120_782 0 0.008f
r152 net10_M1_1120_782 net10_M1_1120_792 1.0
c304 net10_M1_1120_782 0 0.001f
c305 net10_M1_1120_792 0 0.001f
r153 vinp_M1_1760_132 vinp_M1_1760_212 8.0
c306 vinp_M1_1760_132 0 0.008f
c307 vinp_M1_1760_212 0 0.008f
r154 vinp_M1_1760_212 vinp_M1_1760_292 8.0
c308 vinp_M1_1760_212 0 0.008f
c309 vinp_M1_1760_292 0 0.008f
r155 vinp_M1_1760_292 vinp_M1_1760_372 8.0
c310 vinp_M1_1760_292 0 0.008f
c311 vinp_M1_1760_372 0 0.008f
r156 vinp_M1_1760_372 vinp_M1_1760_420 4.8
c312 vinp_M1_1760_372 0 0.0048000000000000004f
c313 vinp_M1_1760_420 0 0.0048000000000000004f
r157 vinp_M1_1760_168 vinp_M1_1760_248 8.0
c314 vinp_M1_1760_168 0 0.008f
c315 vinp_M1_1760_248 0 0.008f
r158 vinp_M1_1760_248 vinp_M1_1760_328 8.0
c316 vinp_M1_1760_248 0 0.008f
c317 vinp_M1_1760_328 0 0.008f
r159 vinp_M1_1760_328 vinp_M1_1760_408 8.0
c318 vinp_M1_1760_328 0 0.008f
c319 vinp_M1_1760_408 0 0.008f
r160 vinp_M1_1760_408 vinp_M1_1760_488 8.0
c320 vinp_M1_1760_408 0 0.008f
c321 vinp_M1_1760_488 0 0.008f
r161 vinp_M1_1760_488 vinp_M1_1760_568 8.0
c322 vinp_M1_1760_488 0 0.008f
c323 vinp_M1_1760_568 0 0.008f
r162 vinp_M1_1760_568 vinp_M1_1760_648 8.0
c324 vinp_M1_1760_568 0 0.008f
c325 vinp_M1_1760_648 0 0.008f
r163 vinp_M1_1760_648 vinp_M1_1760_728 8.0
c326 vinp_M1_1760_648 0 0.008f
c327 vinp_M1_1760_728 0 0.008f
r164 vinp_M1_1760_728 vinp_M1_1760_792 6.4
c328 vinp_M1_1760_728 0 0.0064f
c329 vinp_M1_1760_792 0 0.0064f
r165 net10_M1_1680_132 net10_M1_1680_168 3.5999999999999996
c330 net10_M1_1680_132 0 0.0036f
c331 net10_M1_1680_168 0 0.0036f
r166 net10_M1_1680_168 net10_M1_1680_248 8.0
c332 net10_M1_1680_168 0 0.008f
c333 net10_M1_1680_248 0 0.008f
r167 net10_M1_1680_248 net10_M1_1680_328 8.0
c334 net10_M1_1680_248 0 0.008f
c335 net10_M1_1680_328 0 0.008f
r168 net10_M1_1680_328 net10_M1_1680_336 0.8
c336 net10_M1_1680_328 0 0.0008f
c337 net10_M1_1680_336 0 0.0008f
r169 net10_M1_1680_336 net10_M1_1680_416 8.0
c338 net10_M1_1680_336 0 0.008f
c339 net10_M1_1680_416 0 0.008f
r170 net10_M1_1680_416 net10_M1_1680_462 4.6
c340 net10_M1_1680_416 0 0.0046f
c341 net10_M1_1680_462 0 0.0046f
r171 net10_M1_1680_462 net10_M1_1680_542 8.0
c342 net10_M1_1680_462 0 0.008f
c343 net10_M1_1680_542 0 0.008f
r172 net10_M1_1680_542 net10_M1_1680_588 4.6
c344 net10_M1_1680_542 0 0.0046f
c345 net10_M1_1680_588 0 0.0046f
r173 net10_M1_1680_588 net10_M1_1680_668 8.0
c346 net10_M1_1680_588 0 0.008f
c347 net10_M1_1680_668 0 0.008f
r174 net10_M1_1680_668 net10_M1_1680_748 8.0
c348 net10_M1_1680_668 0 0.008f
c349 net10_M1_1680_748 0 0.008f
r175 net10_M1_1680_748 net10_M1_1680_792 4.3999999999999995
c350 net10_M1_1680_748 0 0.0044f
c351 net10_M1_1680_792 0 0.0044f
r176 net8_M1_1840_132 net8_M1_1840_212 8.0
c352 net8_M1_1840_132 0 0.008f
c353 net8_M1_1840_212 0 0.008f
r177 net8_M1_1840_212 net8_M1_1840_252 4.0
c354 net8_M1_1840_212 0 0.004f
c355 net8_M1_1840_252 0 0.004f
r178 net8_M1_1840_252 net8_M1_1840_332 8.0
c356 net8_M1_1840_252 0 0.008f
c357 net8_M1_1840_332 0 0.008f
r179 net8_M1_1840_332 net8_M1_1840_336 0.4
c358 net8_M1_1840_332 0 0.0004f
c359 net8_M1_1840_336 0 0.0004f
r180 net8_M1_1840_336 net8_M1_1840_416 8.0
c360 net8_M1_1840_336 0 0.008f
c361 net8_M1_1840_416 0 0.008f
r181 net8_M1_1840_416 net8_M1_1840_462 4.6
c362 net8_M1_1840_416 0 0.0046f
c363 net8_M1_1840_462 0 0.0046f
r182 net8_M1_1840_462 net8_M1_1840_542 8.0
c364 net8_M1_1840_462 0 0.008f
c365 net8_M1_1840_542 0 0.008f
r183 net8_M1_1840_542 net8_M1_1840_588 4.6
c366 net8_M1_1840_542 0 0.0046f
c367 net8_M1_1840_588 0 0.0046f
r184 net8_M1_1840_588 net8_M1_1840_668 8.0
c368 net8_M1_1840_588 0 0.008f
c369 net8_M1_1840_668 0 0.008f
r185 net8_M1_1840_668 net8_M1_1840_748 8.0
c370 net8_M1_1840_668 0 0.008f
c371 net8_M1_1840_748 0 0.008f
r186 net8_M1_1840_748 net8_M1_1840_792 4.3999999999999995
c372 net8_M1_1840_748 0 0.0044f
c373 net8_M1_1840_792 0 0.0044f
r187 vinn_M1_2400_132 vinn_M1_2400_212 8.0
c374 vinn_M1_2400_132 0 0.008f
c375 vinn_M1_2400_212 0 0.008f
r188 vinn_M1_2400_212 vinn_M1_2400_292 8.0
c376 vinn_M1_2400_212 0 0.008f
c377 vinn_M1_2400_292 0 0.008f
r189 vinn_M1_2400_292 vinn_M1_2400_372 8.0
c378 vinn_M1_2400_292 0 0.008f
c379 vinn_M1_2400_372 0 0.008f
r190 vinn_M1_2400_372 vinn_M1_2400_452 8.0
c380 vinn_M1_2400_372 0 0.008f
c381 vinn_M1_2400_452 0 0.008f
r191 vinn_M1_2400_452 vinn_M1_2400_504 5.2
c382 vinn_M1_2400_452 0 0.0052f
c383 vinn_M1_2400_504 0 0.0052f
r192 vinn_M1_2400_168 vinn_M1_2400_248 8.0
c384 vinn_M1_2400_168 0 0.008f
c385 vinn_M1_2400_248 0 0.008f
r193 vinn_M1_2400_248 vinn_M1_2400_328 8.0
c386 vinn_M1_2400_248 0 0.008f
c387 vinn_M1_2400_328 0 0.008f
r194 vinn_M1_2400_328 vinn_M1_2400_408 8.0
c388 vinn_M1_2400_328 0 0.008f
c389 vinn_M1_2400_408 0 0.008f
r195 vinn_M1_2400_408 vinn_M1_2400_488 8.0
c390 vinn_M1_2400_408 0 0.008f
c391 vinn_M1_2400_488 0 0.008f
r196 vinn_M1_2400_488 vinn_M1_2400_568 8.0
c392 vinn_M1_2400_488 0 0.008f
c393 vinn_M1_2400_568 0 0.008f
r197 vinn_M1_2400_568 vinn_M1_2400_648 8.0
c394 vinn_M1_2400_568 0 0.008f
c395 vinn_M1_2400_648 0 0.008f
r198 vinn_M1_2400_648 vinn_M1_2400_728 8.0
c396 vinn_M1_2400_648 0 0.008f
c397 vinn_M1_2400_728 0 0.008f
r199 vinn_M1_2400_728 vinn_M1_2400_792 6.4
c398 vinn_M1_2400_728 0 0.0064f
c399 vinn_M1_2400_792 0 0.0064f
r200 net10_M1_2320_132 net10_M1_2320_168 3.5999999999999996
c400 net10_M1_2320_132 0 0.0036f
c401 net10_M1_2320_168 0 0.0036f
r201 net10_M1_2320_168 net10_M1_2320_248 8.0
c402 net10_M1_2320_168 0 0.008f
c403 net10_M1_2320_248 0 0.008f
r202 net10_M1_2320_248 net10_M1_2320_328 8.0
c404 net10_M1_2320_248 0 0.008f
c405 net10_M1_2320_328 0 0.008f
r203 net10_M1_2320_328 net10_M1_2320_336 0.8
c406 net10_M1_2320_328 0 0.0008f
c407 net10_M1_2320_336 0 0.0008f
r204 net10_M1_2320_336 net10_M1_2320_416 8.0
c408 net10_M1_2320_336 0 0.008f
c409 net10_M1_2320_416 0 0.008f
r205 net10_M1_2320_416 net10_M1_2320_462 4.6
c410 net10_M1_2320_416 0 0.0046f
c411 net10_M1_2320_462 0 0.0046f
r206 net10_M1_2320_462 net10_M1_2320_542 8.0
c412 net10_M1_2320_462 0 0.008f
c413 net10_M1_2320_542 0 0.008f
r207 net10_M1_2320_542 net10_M1_2320_588 4.6
c414 net10_M1_2320_542 0 0.0046f
c415 net10_M1_2320_588 0 0.0046f
r208 net10_M1_2320_588 net10_M1_2320_668 8.0
c416 net10_M1_2320_588 0 0.008f
c417 net10_M1_2320_668 0 0.008f
r209 net10_M1_2320_668 net10_M1_2320_748 8.0
c418 net10_M1_2320_668 0 0.008f
c419 net10_M1_2320_748 0 0.008f
r210 net10_M1_2320_748 net10_M1_2320_792 4.3999999999999995
c420 net10_M1_2320_748 0 0.0044f
c421 net10_M1_2320_792 0 0.0044f
r211 vout_M1_2480_132 vout_M1_2480_212 8.0
c422 vout_M1_2480_132 0 0.008f
c423 vout_M1_2480_212 0 0.008f
r212 vout_M1_2480_212 vout_M1_2480_292 8.0
c424 vout_M1_2480_212 0 0.008f
c425 vout_M1_2480_292 0 0.008f
r213 vout_M1_2480_292 vout_M1_2480_336 4.3999999999999995
c426 vout_M1_2480_292 0 0.0044f
c427 vout_M1_2480_336 0 0.0044f
r214 vout_M1_2480_336 vout_M1_2480_416 8.0
c428 vout_M1_2480_336 0 0.008f
c429 vout_M1_2480_416 0 0.008f
r215 vout_M1_2480_416 vout_M1_2480_462 4.6
c430 vout_M1_2480_416 0 0.0046f
c431 vout_M1_2480_462 0 0.0046f
r216 vout_M1_2480_462 vout_M1_2480_542 8.0
c432 vout_M1_2480_462 0 0.008f
c433 vout_M1_2480_542 0 0.008f
r217 vout_M1_2480_542 vout_M1_2480_588 4.6
c434 vout_M1_2480_542 0 0.0046f
c435 vout_M1_2480_588 0 0.0046f
r218 vout_M1_2480_588 vout_M1_2480_668 8.0
c436 vout_M1_2480_588 0 0.008f
c437 vout_M1_2480_668 0 0.008f
r219 vout_M1_2480_668 vout_M1_2480_748 8.0
c438 vout_M1_2480_668 0 0.008f
c439 vout_M1_2480_748 0 0.008f
r220 vout_M1_2480_748 vout_M1_2480_792 4.3999999999999995
c440 vout_M1_2480_748 0 0.0044f
c441 vout_M1_2480_792 0 0.0044f
r221 vss_M2_284_168 vss_M2_364_168 4.8
c442 vss_M2_284_168 0 0.008f
c443 vss_M2_364_168 0 0.008f
r222 vss_M2_364_168 vss_M2_444_168 4.8
c444 vss_M2_364_168 0 0.008f
c445 vss_M2_444_168 0 0.008f
r223 vss_M2_444_168 vss_M2_524_168 4.8
c446 vss_M2_444_168 0 0.008f
c447 vss_M2_524_168 0 0.008f
r224 vss_M2_524_168 vss_M2_604_168 4.8
c448 vss_M2_524_168 0 0.008f
c449 vss_M2_604_168 0 0.008f
r225 vss_M2_604_168 vss_M2_684_168 4.8
c450 vss_M2_604_168 0 0.008f
c451 vss_M2_684_168 0 0.008f
r226 vss_M2_684_168 vss_M2_764_168 4.8
c452 vss_M2_684_168 0 0.008f
c453 vss_M2_764_168 0 0.008f
r227 vss_M2_764_168 vss_M2_844_168 4.8
c454 vss_M2_764_168 0 0.008f
c455 vss_M2_844_168 0 0.008f
r228 vss_M2_844_168 vss_M2_924_168 4.8
c456 vss_M2_844_168 0 0.008f
c457 vss_M2_924_168 0 0.008f
r229 vss_M2_924_168 vss_M2_1004_168 4.8
c458 vss_M2_924_168 0 0.008f
c459 vss_M2_1004_168 0 0.008f
r230 vss_M2_1004_168 vss_M2_1084_168 4.8
c460 vss_M2_1004_168 0 0.008f
c461 vss_M2_1084_168 0 0.008f
r231 vss_M2_1084_168 vss_M2_1164_168 4.8
c462 vss_M2_1084_168 0 0.008f
c463 vss_M2_1164_168 0 0.008f
r232 vss_M2_1164_168 vss_M2_1244_168 4.8
c464 vss_M2_1164_168 0 0.008f
c465 vss_M2_1244_168 0 0.008f
r233 vss_M2_1244_168 vss_M2_1324_168 4.8
c466 vss_M2_1244_168 0 0.008f
c467 vss_M2_1324_168 0 0.008f
r234 vss_M2_1324_168 vss_M2_1404_168 4.8
c468 vss_M2_1324_168 0 0.008f
c469 vss_M2_1404_168 0 0.008f
r235 vss_M2_1404_168 vss_M2_1484_168 4.8
c470 vss_M2_1404_168 0 0.008f
c471 vss_M2_1484_168 0 0.008f
r236 vss_M2_1484_168 vss_M2_1564_168 4.8
c472 vss_M2_1484_168 0 0.008f
c473 vss_M2_1564_168 0 0.008f
r237 vss_M2_1564_168 vss_M2_1644_168 4.8
c474 vss_M2_1564_168 0 0.008f
c475 vss_M2_1644_168 0 0.008f
r238 vss_M2_1644_168 vss_M2_1724_168 4.8
c476 vss_M2_1644_168 0 0.008f
c477 vss_M2_1724_168 0 0.008f
r239 vss_M2_1724_168 vss_M2_1804_168 4.8
c478 vss_M2_1724_168 0 0.008f
c479 vss_M2_1804_168 0 0.008f
r240 vss_M2_1804_168 vss_M2_1884_168 4.8
c480 vss_M2_1804_168 0 0.008f
c481 vss_M2_1884_168 0 0.008f
r241 vss_M2_1884_168 vss_M2_1964_168 4.8
c482 vss_M2_1884_168 0 0.008f
c483 vss_M2_1964_168 0 0.008f
r242 vss_M2_1964_168 vss_M2_2044_168 4.8
c484 vss_M2_1964_168 0 0.008f
c485 vss_M2_2044_168 0 0.008f
r243 vss_M2_2044_168 vss_M2_2124_168 4.8
c486 vss_M2_2044_168 0 0.008f
c487 vss_M2_2124_168 0 0.008f
r244 vss_M2_2124_168 vss_M2_2204_168 4.8
c488 vss_M2_2124_168 0 0.008f
c489 vss_M2_2204_168 0 0.008f
r245 vss_M2_2204_168 vss_M2_2284_168 4.8
c490 vss_M2_2204_168 0 0.008f
c491 vss_M2_2284_168 0 0.008f
r246 vss_M2_2284_168 vss_M2_2364_168 4.8
c492 vss_M2_2284_168 0 0.008f
c493 vss_M2_2364_168 0 0.008f
r247 vss_M2_2364_168 vss_M2_2444_168 4.8
c494 vss_M2_2364_168 0 0.008f
c495 vss_M2_2444_168 0 0.008f
r248 vss_M2_2444_168 vss_M2_2524_168 4.8
c496 vss_M2_2444_168 0 0.008f
c497 vss_M2_2524_168 0 0.008f
r249 vss_M2_2524_168 vss_M2_2604_168 4.8
c498 vss_M2_2524_168 0 0.008f
c499 vss_M2_2604_168 0 0.008f
r250 vss_M2_2604_168 vss_M2_2684_168 4.8
c500 vss_M2_2604_168 0 0.008f
c501 vss_M2_2684_168 0 0.008f
r251 vss_M2_2684_168 vss_M2_2764_168 4.8
c502 vss_M2_2684_168 0 0.008f
c503 vss_M2_2764_168 0 0.008f
r252 vss_M2_2764_168 vss_M2_2844_168 4.8
c504 vss_M2_2764_168 0 0.008f
c505 vss_M2_2844_168 0 0.008f
r253 vss_M2_2844_168 vss_M2_2924_168 4.8
c506 vss_M2_2844_168 0 0.008f
c507 vss_M2_2924_168 0 0.008f
r254 vss_M2_2924_168 vss_M2_3004_168 4.8
c508 vss_M2_2924_168 0 0.008f
c509 vss_M2_3004_168 0 0.008f
r255 vss_M2_3004_168 vss_M2_3084_168 4.8
c510 vss_M2_3004_168 0 0.008f
c511 vss_M2_3084_168 0 0.008f
r256 vss_M2_3084_168 vss_M2_3164_168 4.8
c512 vss_M2_3084_168 0 0.008f
c513 vss_M2_3164_168 0 0.008f
r257 vss_M2_3164_168 vss_M2_3244_168 4.8
c514 vss_M2_3164_168 0 0.008f
c515 vss_M2_3244_168 0 0.008f
r258 vss_M2_3244_168 vss_M2_3324_168 4.8
c516 vss_M2_3244_168 0 0.008f
c517 vss_M2_3324_168 0 0.008f
r259 vss_M2_3324_168 vss_M2_3404_168 4.8
c518 vss_M2_3324_168 0 0.008f
c519 vss_M2_3404_168 0 0.008f
r260 vss_M2_3404_168 vss_M2_3484_168 4.8
c520 vss_M2_3404_168 0 0.008f
c521 vss_M2_3484_168 0 0.008f
r261 vss_M2_3484_168 vss_M2_3564_168 4.8
c522 vss_M2_3484_168 0 0.008f
c523 vss_M2_3564_168 0 0.008f
r262 vss_M2_3564_168 vss_M2_3644_168 4.8
c524 vss_M2_3564_168 0 0.008f
c525 vss_M2_3644_168 0 0.008f
r263 vss_M2_3644_168 vss_M2_3724_168 4.8
c526 vss_M2_3644_168 0 0.008f
c527 vss_M2_3724_168 0 0.008f
r264 vss_M2_3724_168 vss_M2_3804_168 4.8
c528 vss_M2_3724_168 0 0.008f
c529 vss_M2_3804_168 0 0.008f
r265 vss_M2_3804_168 vss_M2_3884_168 4.8
c530 vss_M2_3804_168 0 0.008f
c531 vss_M2_3884_168 0 0.008f
r266 vss_M2_3884_168 vss_M2_3920_168 2.1599999999999997
c532 vss_M2_3884_168 0 0.0036f
c533 vss_M2_3920_168 0 0.0036f
r267 net10_M2_1244_168 net10_M2_1324_168 4.8
c534 net10_M2_1244_168 0 0.008f
c535 net10_M2_1324_168 0 0.008f
r268 net10_M2_1324_168 net10_M2_1404_168 4.8
c536 net10_M2_1324_168 0 0.008f
c537 net10_M2_1404_168 0 0.008f
r269 net10_M2_1404_168 net10_M2_1484_168 4.8
c538 net10_M2_1404_168 0 0.008f
c539 net10_M2_1484_168 0 0.008f
r270 net10_M2_1484_168 net10_M2_1564_168 4.8
c540 net10_M2_1484_168 0 0.008f
c541 net10_M2_1564_168 0 0.008f
r271 net10_M2_1564_168 net10_M2_1644_168 4.8
c542 net10_M2_1564_168 0 0.008f
c543 net10_M2_1644_168 0 0.008f
r272 net10_M2_1644_168 net10_M2_1724_168 4.8
c544 net10_M2_1644_168 0 0.008f
c545 net10_M2_1724_168 0 0.008f
r273 net10_M2_1724_168 net10_M2_1804_168 4.8
c546 net10_M2_1724_168 0 0.008f
c547 net10_M2_1804_168 0 0.008f
r274 net10_M2_1804_168 net10_M2_1884_168 4.8
c548 net10_M2_1804_168 0 0.008f
c549 net10_M2_1884_168 0 0.008f
r275 net10_M2_1884_168 net10_M2_1964_168 4.8
c550 net10_M2_1884_168 0 0.008f
c551 net10_M2_1964_168 0 0.008f
r276 net10_M2_1964_168 net10_M2_2044_168 4.8
c552 net10_M2_1964_168 0 0.008f
c553 net10_M2_2044_168 0 0.008f
r277 net10_M2_2044_168 net10_M2_2124_168 4.8
c554 net10_M2_2044_168 0 0.008f
c555 net10_M2_2124_168 0 0.008f
r278 net10_M2_2124_168 net10_M2_2204_168 4.8
c556 net10_M2_2124_168 0 0.008f
c557 net10_M2_2204_168 0 0.008f
r279 net10_M2_2204_168 net10_M2_2284_168 4.8
c558 net10_M2_2204_168 0 0.008f
c559 net10_M2_2284_168 0 0.008f
r280 net10_M2_2284_168 net10_M2_2364_168 4.8
c560 net10_M2_2284_168 0 0.008f
c561 net10_M2_2364_168 0 0.008f
r281 net10_M2_2364_168 net10_M2_2444_168 4.8
c562 net10_M2_2364_168 0 0.008f
c563 net10_M2_2444_168 0 0.008f
r282 net10_M2_2444_168 net10_M2_2524_168 4.8
c564 net10_M2_2444_168 0 0.008f
c565 net10_M2_2524_168 0 0.008f
r283 net10_M2_2524_168 net10_M2_2604_168 4.8
c566 net10_M2_2524_168 0 0.008f
c567 net10_M2_2604_168 0 0.008f
r284 net10_M2_2604_168 net10_M2_2684_168 4.8
c568 net10_M2_2604_168 0 0.008f
c569 net10_M2_2684_168 0 0.008f
r285 net10_M2_2684_168 net10_M2_2764_168 4.8
c570 net10_M2_2684_168 0 0.008f
c571 net10_M2_2764_168 0 0.008f
r286 net10_M2_2764_168 net10_M2_2844_168 4.8
c572 net10_M2_2764_168 0 0.008f
c573 net10_M2_2844_168 0 0.008f
r287 net10_M2_2844_168 net10_M2_2924_168 4.8
c574 net10_M2_2844_168 0 0.008f
c575 net10_M2_2924_168 0 0.008f
r288 net10_M2_2924_168 net10_M2_3004_168 4.8
c576 net10_M2_2924_168 0 0.008f
c577 net10_M2_3004_168 0 0.008f
r289 net10_M2_3004_168 net10_M2_3084_168 4.8
c578 net10_M2_3004_168 0 0.008f
c579 net10_M2_3084_168 0 0.008f
r290 net10_M2_3084_168 net10_M2_3164_168 4.8
c580 net10_M2_3084_168 0 0.008f
c581 net10_M2_3164_168 0 0.008f
r291 net10_M2_3164_168 net10_M2_3244_168 4.8
c582 net10_M2_3164_168 0 0.008f
c583 net10_M2_3244_168 0 0.008f
r292 net10_M2_3244_168 net10_M2_3324_168 4.8
c584 net10_M2_3244_168 0 0.008f
c585 net10_M2_3324_168 0 0.008f
r293 net10_M2_3324_168 net10_M2_3404_168 4.8
c586 net10_M2_3324_168 0 0.008f
c587 net10_M2_3404_168 0 0.008f
r294 net10_M2_3404_168 net10_M2_3484_168 4.8
c588 net10_M2_3404_168 0 0.008f
c589 net10_M2_3484_168 0 0.008f
r295 net10_M2_3484_168 net10_M2_3564_168 4.8
c590 net10_M2_3484_168 0 0.008f
c591 net10_M2_3564_168 0 0.008f
r296 net10_M2_3564_168 net10_M2_3644_168 4.8
c592 net10_M2_3564_168 0 0.008f
c593 net10_M2_3644_168 0 0.008f
r297 net10_M2_3644_168 net10_M2_3724_168 4.8
c594 net10_M2_3644_168 0 0.008f
c595 net10_M2_3724_168 0 0.008f
r298 net10_M2_3724_168 net10_M2_3804_168 4.8
c596 net10_M2_3724_168 0 0.008f
c597 net10_M2_3804_168 0 0.008f
r299 net10_M2_3804_168 net10_M2_3884_168 4.8
c598 net10_M2_3804_168 0 0.008f
c599 net10_M2_3884_168 0 0.008f
r300 net10_M2_3884_168 net10_M2_3920_168 2.1599999999999997
c600 net10_M2_3884_168 0 0.0036f
c601 net10_M2_3920_168 0 0.0036f
r301 vdd_M2_3004_168 vdd_M2_3084_168 4.8
c602 vdd_M2_3004_168 0 0.008f
c603 vdd_M2_3084_168 0 0.008f
r302 vdd_M2_3084_168 vdd_M2_3164_168 4.8
c604 vdd_M2_3084_168 0 0.008f
c605 vdd_M2_3164_168 0 0.008f
r303 vdd_M2_3164_168 vdd_M2_3244_168 4.8
c606 vdd_M2_3164_168 0 0.008f
c607 vdd_M2_3244_168 0 0.008f
r304 vdd_M2_3244_168 vdd_M2_3324_168 4.8
c608 vdd_M2_3244_168 0 0.008f
c609 vdd_M2_3324_168 0 0.008f
r305 vdd_M2_3324_168 vdd_M2_3404_168 4.8
c610 vdd_M2_3324_168 0 0.008f
c611 vdd_M2_3404_168 0 0.008f
r306 vdd_M2_3404_168 vdd_M2_3484_168 4.8
c612 vdd_M2_3404_168 0 0.008f
c613 vdd_M2_3484_168 0 0.008f
r307 vdd_M2_3484_168 vdd_M2_3564_168 4.8
c614 vdd_M2_3484_168 0 0.008f
c615 vdd_M2_3564_168 0 0.008f
r308 vdd_M2_3564_168 vdd_M2_3644_168 4.8
c616 vdd_M2_3564_168 0 0.008f
c617 vdd_M2_3644_168 0 0.008f
r309 vdd_M2_3644_168 vdd_M2_3724_168 4.8
c618 vdd_M2_3644_168 0 0.008f
c619 vdd_M2_3724_168 0 0.008f
r310 vdd_M2_3724_168 vdd_M2_3804_168 4.8
c620 vdd_M2_3724_168 0 0.008f
c621 vdd_M2_3804_168 0 0.008f
r311 vdd_M2_3804_168 vdd_M2_3884_168 4.8
c622 vdd_M2_3804_168 0 0.008f
c623 vdd_M2_3884_168 0 0.008f
r312 vdd_M2_3884_168 vdd_M2_3920_168 2.1599999999999997
c624 vdd_M2_3884_168 0 0.0036f
c625 vdd_M2_3920_168 0 0.0036f
r313 vdd_M2_320_168 vdd_M2_400_168 4.8
c626 vdd_M2_320_168 0 0.008f
c627 vdd_M2_400_168 0 0.008f
r314 vdd_M2_400_168 vdd_M2_480_168 4.8
c628 vdd_M2_400_168 0 0.008f
c629 vdd_M2_480_168 0 0.008f
r315 vdd_M2_480_168 vdd_M2_560_168 4.8
c630 vdd_M2_480_168 0 0.008f
c631 vdd_M2_560_168 0 0.008f
r316 vdd_M2_560_168 vdd_M2_640_168 4.8
c632 vdd_M2_560_168 0 0.008f
c633 vdd_M2_640_168 0 0.008f
r317 vdd_M2_640_168 vdd_M2_720_168 4.8
c634 vdd_M2_640_168 0 0.008f
c635 vdd_M2_720_168 0 0.008f
r318 vdd_M2_720_168 vdd_M2_800_168 4.8
c636 vdd_M2_720_168 0 0.008f
c637 vdd_M2_800_168 0 0.008f
r319 vdd_M2_800_168 vdd_M2_880_168 4.8
c638 vdd_M2_800_168 0 0.008f
c639 vdd_M2_880_168 0 0.008f
r320 vdd_M2_880_168 vdd_M2_960_168 4.8
c640 vdd_M2_880_168 0 0.008f
c641 vdd_M2_960_168 0 0.008f
r321 vdd_M2_960_168 vdd_M2_1040_168 4.8
c642 vdd_M2_960_168 0 0.008f
c643 vdd_M2_1040_168 0 0.008f
r322 vdd_M2_1040_168 vdd_M2_1120_168 4.8
c644 vdd_M2_1040_168 0 0.008f
c645 vdd_M2_1120_168 0 0.008f
r323 vdd_M2_1120_168 vdd_M2_1200_168 4.8
c646 vdd_M2_1120_168 0 0.008f
c647 vdd_M2_1200_168 0 0.008f
r324 vdd_M2_1200_168 vdd_M2_1280_168 4.8
c648 vdd_M2_1200_168 0 0.008f
c649 vdd_M2_1280_168 0 0.008f
r325 vdd_M2_1280_168 vdd_M2_1360_168 4.8
c650 vdd_M2_1280_168 0 0.008f
c651 vdd_M2_1360_168 0 0.008f
r326 vdd_M2_1360_168 vdd_M2_1440_168 4.8
c652 vdd_M2_1360_168 0 0.008f
c653 vdd_M2_1440_168 0 0.008f
r327 vdd_M2_1440_168 vdd_M2_1520_168 4.8
c654 vdd_M2_1440_168 0 0.008f
c655 vdd_M2_1520_168 0 0.008f
r328 vdd_M2_1520_168 vdd_M2_1600_168 4.8
c656 vdd_M2_1520_168 0 0.008f
c657 vdd_M2_1600_168 0 0.008f
r329 vdd_M2_1600_168 vdd_M2_1680_168 4.8
c658 vdd_M2_1600_168 0 0.008f
c659 vdd_M2_1680_168 0 0.008f
r330 vdd_M2_1680_168 vdd_M2_1760_168 4.8
c660 vdd_M2_1680_168 0 0.008f
c661 vdd_M2_1760_168 0 0.008f
r331 vdd_M2_1760_168 vdd_M2_1840_168 4.8
c662 vdd_M2_1760_168 0 0.008f
c663 vdd_M2_1840_168 0 0.008f
r332 vdd_M2_1840_168 vdd_M2_1920_168 4.8
c664 vdd_M2_1840_168 0 0.008f
c665 vdd_M2_1920_168 0 0.008f
r333 vdd_M2_1920_168 vdd_M2_2000_168 4.8
c666 vdd_M2_1920_168 0 0.008f
c667 vdd_M2_2000_168 0 0.008f
r334 vdd_M2_2000_168 vdd_M2_2080_168 4.8
c668 vdd_M2_2000_168 0 0.008f
c669 vdd_M2_2080_168 0 0.008f
r335 vdd_M2_2080_168 vdd_M2_2160_168 4.8
c670 vdd_M2_2080_168 0 0.008f
c671 vdd_M2_2160_168 0 0.008f
r336 vdd_M2_2160_168 vdd_M2_2240_168 4.8
c672 vdd_M2_2160_168 0 0.008f
c673 vdd_M2_2240_168 0 0.008f
r337 vdd_M2_2240_168 vdd_M2_2320_168 4.8
c674 vdd_M2_2240_168 0 0.008f
c675 vdd_M2_2320_168 0 0.008f
r338 vdd_M2_2320_168 vdd_M2_2400_168 4.8
c676 vdd_M2_2320_168 0 0.008f
c677 vdd_M2_2400_168 0 0.008f
r339 vdd_M2_2400_168 vdd_M2_2480_168 4.8
c678 vdd_M2_2400_168 0 0.008f
c679 vdd_M2_2480_168 0 0.008f
r340 vdd_M2_2480_168 vdd_M2_2560_168 4.8
c680 vdd_M2_2480_168 0 0.008f
c681 vdd_M2_2560_168 0 0.008f
r341 vdd_M2_2560_168 vdd_M2_2640_168 4.8
c682 vdd_M2_2560_168 0 0.008f
c683 vdd_M2_2640_168 0 0.008f
r342 vdd_M2_2640_168 vdd_M2_2720_168 4.8
c684 vdd_M2_2640_168 0 0.008f
c685 vdd_M2_2720_168 0 0.008f
r343 vdd_M2_2720_168 vdd_M2_2800_168 4.8
c686 vdd_M2_2720_168 0 0.008f
c687 vdd_M2_2800_168 0 0.008f
r344 vdd_M2_2800_168 vdd_M2_2880_168 4.8
c688 vdd_M2_2800_168 0 0.008f
c689 vdd_M2_2880_168 0 0.008f
r345 vdd_M2_2880_168 vdd_M2_2960_168 4.8
c690 vdd_M2_2880_168 0 0.008f
c691 vdd_M2_2960_168 0 0.008f
r346 vdd_M2_2960_168 vdd_M2_3040_168 4.8
c692 vdd_M2_2960_168 0 0.008f
c693 vdd_M2_3040_168 0 0.008f
r347 vdd_M2_3040_168 vdd_M2_3120_168 4.8
c694 vdd_M2_3040_168 0 0.008f
c695 vdd_M2_3120_168 0 0.008f
r348 vdd_M2_3120_168 vdd_M2_3200_168 4.8
c696 vdd_M2_3120_168 0 0.008f
c697 vdd_M2_3200_168 0 0.008f
r349 vdd_M2_3200_168 vdd_M2_3280_168 4.8
c698 vdd_M2_3200_168 0 0.008f
c699 vdd_M2_3280_168 0 0.008f
r350 vdd_M2_3280_168 vdd_M2_3316_168 2.1599999999999997
c700 vdd_M2_3280_168 0 0.0036f
c701 vdd_M2_3316_168 0 0.0036f
r351 vdd_M2_3280_168 vdd_M2_3360_168 4.8
c702 vdd_M2_3280_168 0 0.008f
c703 vdd_M2_3360_168 0 0.008f
r352 vdd_M2_3360_168 vdd_M2_3440_168 4.8
c704 vdd_M2_3360_168 0 0.008f
c705 vdd_M2_3440_168 0 0.008f
r353 vdd_M2_3440_168 vdd_M2_3520_168 4.8
c706 vdd_M2_3440_168 0 0.008f
c707 vdd_M2_3520_168 0 0.008f
r354 vdd_M2_3520_168 vdd_M2_3600_168 4.8
c708 vdd_M2_3520_168 0 0.008f
c709 vdd_M2_3600_168 0 0.008f
r355 vdd_M2_3600_168 vdd_M2_3680_168 4.8
c710 vdd_M2_3600_168 0 0.008f
c711 vdd_M2_3680_168 0 0.008f
r356 vdd_M2_3680_168 vdd_M2_3760_168 4.8
c712 vdd_M2_3680_168 0 0.008f
c713 vdd_M2_3760_168 0 0.008f
r357 vdd_M2_3760_168 vdd_M2_3840_168 4.8
c714 vdd_M2_3760_168 0 0.008f
c715 vdd_M2_3840_168 0 0.008f
r358 vdd_M2_3840_168 vdd_M2_3920_168 4.8
c716 vdd_M2_3840_168 0 0.008f
c717 vdd_M2_3920_168 0 0.008f
r359 vdd_M2_3920_168 vdd_M2_3956_168 2.1599999999999997
c718 vdd_M2_3920_168 0 0.0036f
c719 vdd_M2_3956_168 0 0.0036f
r360 net10_M2_684_336 net10_M2_764_336 4.8
c720 net10_M2_684_336 0 0.008f
c721 net10_M2_764_336 0 0.008f
r361 net10_M2_764_336 net10_M2_844_336 4.8
c722 net10_M2_764_336 0 0.008f
c723 net10_M2_844_336 0 0.008f
r362 net10_M2_844_336 net10_M2_924_336 4.8
c724 net10_M2_844_336 0 0.008f
c725 net10_M2_924_336 0 0.008f
r363 net10_M2_924_336 net10_M2_1004_336 4.8
c726 net10_M2_924_336 0 0.008f
c727 net10_M2_1004_336 0 0.008f
r364 net10_M2_1004_336 net10_M2_1084_336 4.8
c728 net10_M2_1004_336 0 0.008f
c729 net10_M2_1084_336 0 0.008f
r365 net10_M2_1084_336 net10_M2_1164_336 4.8
c730 net10_M2_1084_336 0 0.008f
c731 net10_M2_1164_336 0 0.008f
r366 net10_M2_1164_336 net10_M2_1244_336 4.8
c732 net10_M2_1164_336 0 0.008f
c733 net10_M2_1244_336 0 0.008f
r367 net10_M2_1244_336 net10_M2_1324_336 4.8
c734 net10_M2_1244_336 0 0.008f
c735 net10_M2_1324_336 0 0.008f
r368 net10_M2_1324_336 net10_M2_1404_336 4.8
c736 net10_M2_1324_336 0 0.008f
c737 net10_M2_1404_336 0 0.008f
r369 net10_M2_1404_336 net10_M2_1484_336 4.8
c738 net10_M2_1404_336 0 0.008f
c739 net10_M2_1484_336 0 0.008f
r370 net10_M2_1484_336 net10_M2_1564_336 4.8
c740 net10_M2_1484_336 0 0.008f
c741 net10_M2_1564_336 0 0.008f
r371 net10_M2_1564_336 net10_M2_1644_336 4.8
c742 net10_M2_1564_336 0 0.008f
c743 net10_M2_1644_336 0 0.008f
r372 net10_M2_1644_336 net10_M2_1724_336 4.8
c744 net10_M2_1644_336 0 0.008f
c745 net10_M2_1724_336 0 0.008f
r373 net10_M2_1724_336 net10_M2_1804_336 4.8
c746 net10_M2_1724_336 0 0.008f
c747 net10_M2_1804_336 0 0.008f
r374 net10_M2_1804_336 net10_M2_1884_336 4.8
c748 net10_M2_1804_336 0 0.008f
c749 net10_M2_1884_336 0 0.008f
r375 net10_M2_1884_336 net10_M2_1964_336 4.8
c750 net10_M2_1884_336 0 0.008f
c751 net10_M2_1964_336 0 0.008f
r376 net10_M2_1964_336 net10_M2_2044_336 4.8
c752 net10_M2_1964_336 0 0.008f
c753 net10_M2_2044_336 0 0.008f
r377 net10_M2_2044_336 net10_M2_2124_336 4.8
c754 net10_M2_2044_336 0 0.008f
c755 net10_M2_2124_336 0 0.008f
r378 net10_M2_2124_336 net10_M2_2204_336 4.8
c756 net10_M2_2124_336 0 0.008f
c757 net10_M2_2204_336 0 0.008f
r379 net10_M2_2204_336 net10_M2_2284_336 4.8
c758 net10_M2_2204_336 0 0.008f
c759 net10_M2_2284_336 0 0.008f
r380 net10_M2_2284_336 net10_M2_2364_336 4.8
c760 net10_M2_2284_336 0 0.008f
c761 net10_M2_2364_336 0 0.008f
r381 net10_M2_2364_336 net10_M2_2444_336 4.8
c762 net10_M2_2364_336 0 0.008f
c763 net10_M2_2444_336 0 0.008f
r382 net10_M2_2444_336 net10_M2_2524_336 4.8
c764 net10_M2_2444_336 0 0.008f
c765 net10_M2_2524_336 0 0.008f
r383 net10_M2_2524_336 net10_M2_2604_336 4.8
c766 net10_M2_2524_336 0 0.008f
c767 net10_M2_2604_336 0 0.008f
r384 net10_M2_2604_336 net10_M2_2684_336 4.8
c768 net10_M2_2604_336 0 0.008f
c769 net10_M2_2684_336 0 0.008f
r385 net10_M2_2684_336 net10_M2_2764_336 4.8
c770 net10_M2_2684_336 0 0.008f
c771 net10_M2_2764_336 0 0.008f
r386 net10_M2_2764_336 net10_M2_2844_336 4.8
c772 net10_M2_2764_336 0 0.008f
c773 net10_M2_2844_336 0 0.008f
r387 net10_M2_2844_336 net10_M2_2924_336 4.8
c774 net10_M2_2844_336 0 0.008f
c775 net10_M2_2924_336 0 0.008f
r388 net10_M2_2924_336 net10_M2_3004_336 4.8
c776 net10_M2_2924_336 0 0.008f
c777 net10_M2_3004_336 0 0.008f
r389 net10_M2_3004_336 net10_M2_3084_336 4.8
c778 net10_M2_3004_336 0 0.008f
c779 net10_M2_3084_336 0 0.008f
r390 net10_M2_3084_336 net10_M2_3164_336 4.8
c780 net10_M2_3084_336 0 0.008f
c781 net10_M2_3164_336 0 0.008f
r391 net10_M2_3164_336 net10_M2_3244_336 4.8
c782 net10_M2_3164_336 0 0.008f
c783 net10_M2_3244_336 0 0.008f
r392 net10_M2_3244_336 net10_M2_3324_336 4.8
c784 net10_M2_3244_336 0 0.008f
c785 net10_M2_3324_336 0 0.008f
r393 net10_M2_3324_336 net10_M2_3404_336 4.8
c786 net10_M2_3324_336 0 0.008f
c787 net10_M2_3404_336 0 0.008f
r394 net10_M2_3404_336 net10_M2_3484_336 4.8
c788 net10_M2_3404_336 0 0.008f
c789 net10_M2_3484_336 0 0.008f
r395 net10_M2_3484_336 net10_M2_3564_336 4.8
c790 net10_M2_3484_336 0 0.008f
c791 net10_M2_3564_336 0 0.008f
r396 net10_M2_3564_336 net10_M2_3644_336 4.8
c792 net10_M2_3564_336 0 0.008f
c793 net10_M2_3644_336 0 0.008f
r397 net10_M2_3644_336 net10_M2_3724_336 4.8
c794 net10_M2_3644_336 0 0.008f
c795 net10_M2_3724_336 0 0.008f
r398 net10_M2_3724_336 net10_M2_3804_336 4.8
c796 net10_M2_3724_336 0 0.008f
c797 net10_M2_3804_336 0 0.008f
r399 net10_M2_3804_336 net10_M2_3884_336 4.8
c798 net10_M2_3804_336 0 0.008f
c799 net10_M2_3884_336 0 0.008f
r400 net10_M2_3884_336 net10_M2_3920_336 2.1599999999999997
c800 net10_M2_3884_336 0 0.0036f
c801 net10_M2_3920_336 0 0.0036f
r401 vout_M2_2284_336 vout_M2_2364_336 4.8
c802 vout_M2_2284_336 0 0.008f
c803 vout_M2_2364_336 0 0.008f
r402 vout_M2_2364_336 vout_M2_2444_336 4.8
c804 vout_M2_2364_336 0 0.008f
c805 vout_M2_2444_336 0 0.008f
r403 vout_M2_2444_336 vout_M2_2524_336 4.8
c806 vout_M2_2444_336 0 0.008f
c807 vout_M2_2524_336 0 0.008f
r404 vout_M2_2524_336 vout_M2_2604_336 4.8
c808 vout_M2_2524_336 0 0.008f
c809 vout_M2_2604_336 0 0.008f
r405 vout_M2_2604_336 vout_M2_2684_336 4.8
c810 vout_M2_2604_336 0 0.008f
c811 vout_M2_2684_336 0 0.008f
r406 vout_M2_2684_336 vout_M2_2764_336 4.8
c812 vout_M2_2684_336 0 0.008f
c813 vout_M2_2764_336 0 0.008f
r407 vout_M2_2764_336 vout_M2_2844_336 4.8
c814 vout_M2_2764_336 0 0.008f
c815 vout_M2_2844_336 0 0.008f
r408 vout_M2_2844_336 vout_M2_2924_336 4.8
c816 vout_M2_2844_336 0 0.008f
c817 vout_M2_2924_336 0 0.008f
r409 vout_M2_2924_336 vout_M2_3004_336 4.8
c818 vout_M2_2924_336 0 0.008f
c819 vout_M2_3004_336 0 0.008f
r410 vout_M2_3004_336 vout_M2_3084_336 4.8
c820 vout_M2_3004_336 0 0.008f
c821 vout_M2_3084_336 0 0.008f
r411 vout_M2_3084_336 vout_M2_3164_336 4.8
c822 vout_M2_3084_336 0 0.008f
c823 vout_M2_3164_336 0 0.008f
r412 vout_M2_3164_336 vout_M2_3244_336 4.8
c824 vout_M2_3164_336 0 0.008f
c825 vout_M2_3244_336 0 0.008f
r413 vout_M2_3244_336 vout_M2_3324_336 4.8
c826 vout_M2_3244_336 0 0.008f
c827 vout_M2_3324_336 0 0.008f
r414 vout_M2_3324_336 vout_M2_3404_336 4.8
c828 vout_M2_3324_336 0 0.008f
c829 vout_M2_3404_336 0 0.008f
r415 vout_M2_3404_336 vout_M2_3484_336 4.8
c830 vout_M2_3404_336 0 0.008f
c831 vout_M2_3484_336 0 0.008f
r416 vout_M2_3484_336 vout_M2_3564_336 4.8
c832 vout_M2_3484_336 0 0.008f
c833 vout_M2_3564_336 0 0.008f
r417 vout_M2_3564_336 vout_M2_3644_336 4.8
c834 vout_M2_3564_336 0 0.008f
c835 vout_M2_3644_336 0 0.008f
r418 vout_M2_3644_336 vout_M2_3724_336 4.8
c836 vout_M2_3644_336 0 0.008f
c837 vout_M2_3724_336 0 0.008f
r419 vout_M2_3724_336 vout_M2_3804_336 4.8
c838 vout_M2_3724_336 0 0.008f
c839 vout_M2_3804_336 0 0.008f
r420 vout_M2_3804_336 vout_M2_3884_336 4.8
c840 vout_M2_3804_336 0 0.008f
c841 vout_M2_3884_336 0 0.008f
r421 vout_M2_3884_336 vout_M2_3920_336 2.1599999999999997
c842 vout_M2_3884_336 0 0.0036f
c843 vout_M2_3920_336 0 0.0036f
r422 net8_M2_2844_336 net8_M2_2924_336 4.8
c844 net8_M2_2844_336 0 0.008f
c845 net8_M2_2924_336 0 0.008f
r423 net8_M2_2924_336 net8_M2_3004_336 4.8
c846 net8_M2_2924_336 0 0.008f
c847 net8_M2_3004_336 0 0.008f
r424 net8_M2_3004_336 net8_M2_3084_336 4.8
c848 net8_M2_3004_336 0 0.008f
c849 net8_M2_3084_336 0 0.008f
r425 net8_M2_3084_336 net8_M2_3164_336 4.8
c850 net8_M2_3084_336 0 0.008f
c851 net8_M2_3164_336 0 0.008f
r426 net8_M2_3164_336 net8_M2_3244_336 4.8
c852 net8_M2_3164_336 0 0.008f
c853 net8_M2_3244_336 0 0.008f
r427 net8_M2_3244_336 net8_M2_3324_336 4.8
c854 net8_M2_3244_336 0 0.008f
c855 net8_M2_3324_336 0 0.008f
r428 net8_M2_3324_336 net8_M2_3404_336 4.8
c856 net8_M2_3324_336 0 0.008f
c857 net8_M2_3404_336 0 0.008f
r429 net8_M2_3404_336 net8_M2_3484_336 4.8
c858 net8_M2_3404_336 0 0.008f
c859 net8_M2_3484_336 0 0.008f
r430 net8_M2_3484_336 net8_M2_3564_336 4.8
c860 net8_M2_3484_336 0 0.008f
c861 net8_M2_3564_336 0 0.008f
r431 net8_M2_3564_336 net8_M2_3644_336 4.8
c862 net8_M2_3564_336 0 0.008f
c863 net8_M2_3644_336 0 0.008f
r432 net8_M2_3644_336 net8_M2_3724_336 4.8
c864 net8_M2_3644_336 0 0.008f
c865 net8_M2_3724_336 0 0.008f
r433 net8_M2_3724_336 net8_M2_3804_336 4.8
c866 net8_M2_3724_336 0 0.008f
c867 net8_M2_3804_336 0 0.008f
r434 net8_M2_3804_336 net8_M2_3884_336 4.8
c868 net8_M2_3804_336 0 0.008f
c869 net8_M2_3884_336 0 0.008f
r435 net8_M2_3884_336 net8_M2_3920_336 2.1599999999999997
c870 net8_M2_3884_336 0 0.0036f
c871 net8_M2_3920_336 0 0.0036f
r436 net8_M2_1120_336 net8_M2_1200_336 4.8
c872 net8_M2_1120_336 0 0.008f
c873 net8_M2_1200_336 0 0.008f
r437 net8_M2_1200_336 net8_M2_1280_336 4.8
c874 net8_M2_1200_336 0 0.008f
c875 net8_M2_1280_336 0 0.008f
r438 net8_M2_1280_336 net8_M2_1360_336 4.8
c876 net8_M2_1280_336 0 0.008f
c877 net8_M2_1360_336 0 0.008f
r439 net8_M2_1360_336 net8_M2_1440_336 4.8
c878 net8_M2_1360_336 0 0.008f
c879 net8_M2_1440_336 0 0.008f
r440 net8_M2_1440_336 net8_M2_1520_336 4.8
c880 net8_M2_1440_336 0 0.008f
c881 net8_M2_1520_336 0 0.008f
r441 net8_M2_1520_336 net8_M2_1600_336 4.8
c882 net8_M2_1520_336 0 0.008f
c883 net8_M2_1600_336 0 0.008f
r442 net8_M2_1600_336 net8_M2_1680_336 4.8
c884 net8_M2_1600_336 0 0.008f
c885 net8_M2_1680_336 0 0.008f
r443 net8_M2_1680_336 net8_M2_1760_336 4.8
c886 net8_M2_1680_336 0 0.008f
c887 net8_M2_1760_336 0 0.008f
r444 net8_M2_1760_336 net8_M2_1840_336 4.8
c888 net8_M2_1760_336 0 0.008f
c889 net8_M2_1840_336 0 0.008f
r445 net8_M2_1840_336 net8_M2_1920_336 4.8
c890 net8_M2_1840_336 0 0.008f
c891 net8_M2_1920_336 0 0.008f
r446 net8_M2_1920_336 net8_M2_2000_336 4.8
c892 net8_M2_1920_336 0 0.008f
c893 net8_M2_2000_336 0 0.008f
r447 net8_M2_2000_336 net8_M2_2080_336 4.8
c894 net8_M2_2000_336 0 0.008f
c895 net8_M2_2080_336 0 0.008f
r448 net8_M2_2080_336 net8_M2_2160_336 4.8
c896 net8_M2_2080_336 0 0.008f
c897 net8_M2_2160_336 0 0.008f
r449 net8_M2_2160_336 net8_M2_2240_336 4.8
c898 net8_M2_2160_336 0 0.008f
c899 net8_M2_2240_336 0 0.008f
r450 net8_M2_2240_336 net8_M2_2320_336 4.8
c900 net8_M2_2240_336 0 0.008f
c901 net8_M2_2320_336 0 0.008f
r451 net8_M2_2320_336 net8_M2_2400_336 4.8
c902 net8_M2_2320_336 0 0.008f
c903 net8_M2_2400_336 0 0.008f
r452 net8_M2_2400_336 net8_M2_2480_336 4.8
c904 net8_M2_2400_336 0 0.008f
c905 net8_M2_2480_336 0 0.008f
r453 net8_M2_2480_336 net8_M2_2560_336 4.8
c906 net8_M2_2480_336 0 0.008f
c907 net8_M2_2560_336 0 0.008f
r454 net8_M2_2560_336 net8_M2_2640_336 4.8
c908 net8_M2_2560_336 0 0.008f
c909 net8_M2_2640_336 0 0.008f
r455 net8_M2_2640_336 net8_M2_2720_336 4.8
c910 net8_M2_2640_336 0 0.008f
c911 net8_M2_2720_336 0 0.008f
r456 net8_M2_2720_336 net8_M2_2800_336 4.8
c912 net8_M2_2720_336 0 0.008f
c913 net8_M2_2800_336 0 0.008f
r457 net8_M2_2800_336 net8_M2_2880_336 4.8
c914 net8_M2_2800_336 0 0.008f
c915 net8_M2_2880_336 0 0.008f
r458 net8_M2_2880_336 net8_M2_2960_336 4.8
c916 net8_M2_2880_336 0 0.008f
c917 net8_M2_2960_336 0 0.008f
r459 net8_M2_2960_336 net8_M2_3040_336 4.8
c918 net8_M2_2960_336 0 0.008f
c919 net8_M2_3040_336 0 0.008f
r460 net8_M2_3040_336 net8_M2_3120_336 4.8
c920 net8_M2_3040_336 0 0.008f
c921 net8_M2_3120_336 0 0.008f
r461 net8_M2_3120_336 net8_M2_3200_336 4.8
c922 net8_M2_3120_336 0 0.008f
c923 net8_M2_3200_336 0 0.008f
r462 net8_M2_3200_336 net8_M2_3236_336 2.1599999999999997
c924 net8_M2_3200_336 0 0.0036f
c925 net8_M2_3236_336 0 0.0036f
r463 vdd_M2_3324_336 vdd_M2_3404_336 4.8
c926 vdd_M2_3324_336 0 0.008f
c927 vdd_M2_3404_336 0 0.008f
r464 vdd_M2_3404_336 vdd_M2_3484_336 4.8
c928 vdd_M2_3404_336 0 0.008f
c929 vdd_M2_3484_336 0 0.008f
r465 vdd_M2_3484_336 vdd_M2_3564_336 4.8
c930 vdd_M2_3484_336 0 0.008f
c931 vdd_M2_3564_336 0 0.008f
r466 vdd_M2_3564_336 vdd_M2_3644_336 4.8
c932 vdd_M2_3564_336 0 0.008f
c933 vdd_M2_3644_336 0 0.008f
r467 vdd_M2_3644_336 vdd_M2_3724_336 4.8
c934 vdd_M2_3644_336 0 0.008f
c935 vdd_M2_3724_336 0 0.008f
r468 vdd_M2_3724_336 vdd_M2_3804_336 4.8
c936 vdd_M2_3724_336 0 0.008f
c937 vdd_M2_3804_336 0 0.008f
r469 vdd_M2_3804_336 vdd_M2_3884_336 4.8
c938 vdd_M2_3804_336 0 0.008f
c939 vdd_M2_3884_336 0 0.008f
r470 vdd_M2_3884_336 vdd_M2_3920_336 2.1599999999999997
c940 vdd_M2_3884_336 0 0.0036f
c941 vdd_M2_3920_336 0 0.0036f
r471 vdd_M2_1120_336 vdd_M2_1200_336 4.8
c942 vdd_M2_1120_336 0 0.008f
c943 vdd_M2_1200_336 0 0.008f
r472 vdd_M2_1200_336 vdd_M2_1280_336 4.8
c944 vdd_M2_1200_336 0 0.008f
c945 vdd_M2_1280_336 0 0.008f
r473 vdd_M2_1280_336 vdd_M2_1360_336 4.8
c946 vdd_M2_1280_336 0 0.008f
c947 vdd_M2_1360_336 0 0.008f
r474 vdd_M2_1360_336 vdd_M2_1440_336 4.8
c948 vdd_M2_1360_336 0 0.008f
c949 vdd_M2_1440_336 0 0.008f
r475 vdd_M2_1440_336 vdd_M2_1520_336 4.8
c950 vdd_M2_1440_336 0 0.008f
c951 vdd_M2_1520_336 0 0.008f
r476 vdd_M2_1520_336 vdd_M2_1600_336 4.8
c952 vdd_M2_1520_336 0 0.008f
c953 vdd_M2_1600_336 0 0.008f
r477 vdd_M2_1600_336 vdd_M2_1680_336 4.8
c954 vdd_M2_1600_336 0 0.008f
c955 vdd_M2_1680_336 0 0.008f
r478 vdd_M2_1680_336 vdd_M2_1760_336 4.8
c956 vdd_M2_1680_336 0 0.008f
c957 vdd_M2_1760_336 0 0.008f
r479 vdd_M2_1760_336 vdd_M2_1840_336 4.8
c958 vdd_M2_1760_336 0 0.008f
c959 vdd_M2_1840_336 0 0.008f
r480 vdd_M2_1840_336 vdd_M2_1920_336 4.8
c960 vdd_M2_1840_336 0 0.008f
c961 vdd_M2_1920_336 0 0.008f
r481 vdd_M2_1920_336 vdd_M2_2000_336 4.8
c962 vdd_M2_1920_336 0 0.008f
c963 vdd_M2_2000_336 0 0.008f
r482 vdd_M2_2000_336 vdd_M2_2080_336 4.8
c964 vdd_M2_2000_336 0 0.008f
c965 vdd_M2_2080_336 0 0.008f
r483 vdd_M2_2080_336 vdd_M2_2160_336 4.8
c966 vdd_M2_2080_336 0 0.008f
c967 vdd_M2_2160_336 0 0.008f
r484 vdd_M2_2160_336 vdd_M2_2240_336 4.8
c968 vdd_M2_2160_336 0 0.008f
c969 vdd_M2_2240_336 0 0.008f
r485 vdd_M2_2240_336 vdd_M2_2320_336 4.8
c970 vdd_M2_2240_336 0 0.008f
c971 vdd_M2_2320_336 0 0.008f
r486 vdd_M2_2320_336 vdd_M2_2400_336 4.8
c972 vdd_M2_2320_336 0 0.008f
c973 vdd_M2_2400_336 0 0.008f
r487 vdd_M2_2400_336 vdd_M2_2480_336 4.8
c974 vdd_M2_2400_336 0 0.008f
c975 vdd_M2_2480_336 0 0.008f
r488 vdd_M2_2480_336 vdd_M2_2560_336 4.8
c976 vdd_M2_2480_336 0 0.008f
c977 vdd_M2_2560_336 0 0.008f
r489 vdd_M2_2560_336 vdd_M2_2640_336 4.8
c978 vdd_M2_2560_336 0 0.008f
c979 vdd_M2_2640_336 0 0.008f
r490 vdd_M2_2640_336 vdd_M2_2720_336 4.8
c980 vdd_M2_2640_336 0 0.008f
c981 vdd_M2_2720_336 0 0.008f
r491 vdd_M2_2720_336 vdd_M2_2800_336 4.8
c982 vdd_M2_2720_336 0 0.008f
c983 vdd_M2_2800_336 0 0.008f
r492 vdd_M2_2800_336 vdd_M2_2880_336 4.8
c984 vdd_M2_2800_336 0 0.008f
c985 vdd_M2_2880_336 0 0.008f
r493 vdd_M2_2880_336 vdd_M2_2960_336 4.8
c986 vdd_M2_2880_336 0 0.008f
c987 vdd_M2_2960_336 0 0.008f
r494 vdd_M2_2960_336 vdd_M2_3040_336 4.8
c988 vdd_M2_2960_336 0 0.008f
c989 vdd_M2_3040_336 0 0.008f
r495 vdd_M2_3040_336 vdd_M2_3120_336 4.8
c990 vdd_M2_3040_336 0 0.008f
c991 vdd_M2_3120_336 0 0.008f
r496 vdd_M2_3120_336 vdd_M2_3200_336 4.8
c992 vdd_M2_3120_336 0 0.008f
c993 vdd_M2_3200_336 0 0.008f
r497 vdd_M2_3200_336 vdd_M2_3280_336 4.8
c994 vdd_M2_3200_336 0 0.008f
c995 vdd_M2_3280_336 0 0.008f
r498 vdd_M2_3280_336 vdd_M2_3360_336 4.8
c996 vdd_M2_3280_336 0 0.008f
c997 vdd_M2_3360_336 0 0.008f
r499 vdd_M2_3360_336 vdd_M2_3440_336 4.8
c998 vdd_M2_3360_336 0 0.008f
c999 vdd_M2_3440_336 0 0.008f
r500 vdd_M2_3440_336 vdd_M2_3520_336 4.8
c1000 vdd_M2_3440_336 0 0.008f
c1001 vdd_M2_3520_336 0 0.008f
r501 vdd_M2_3520_336 vdd_M2_3600_336 4.8
c1002 vdd_M2_3520_336 0 0.008f
c1003 vdd_M2_3600_336 0 0.008f
r502 vdd_M2_3600_336 vdd_M2_3636_336 2.1599999999999997
c1004 vdd_M2_3600_336 0 0.0036f
c1005 vdd_M2_3636_336 0 0.0036f
r503 vdd_M2_3600_336 vdd_M2_3680_336 4.8
c1006 vdd_M2_3600_336 0 0.008f
c1007 vdd_M2_3680_336 0 0.008f
r504 vdd_M2_3680_336 vdd_M2_3760_336 4.8
c1008 vdd_M2_3680_336 0 0.008f
c1009 vdd_M2_3760_336 0 0.008f
r505 vdd_M2_720_336 vdd_M2_800_336 4.8
c1010 vdd_M2_720_336 0 0.008f
c1011 vdd_M2_800_336 0 0.008f
r506 vdd_M2_800_336 vdd_M2_880_336 4.8
c1012 vdd_M2_800_336 0 0.008f
c1013 vdd_M2_880_336 0 0.008f
r507 vdd_M2_880_336 vdd_M2_960_336 4.8
c1014 vdd_M2_880_336 0 0.008f
c1015 vdd_M2_960_336 0 0.008f
r508 vdd_M2_960_336 vdd_M2_1040_336 4.8
c1016 vdd_M2_960_336 0 0.008f
c1017 vdd_M2_1040_336 0 0.008f
r509 vdd_M2_1040_336 vdd_M2_1120_336 4.8
c1018 vdd_M2_1040_336 0 0.008f
c1019 vdd_M2_1120_336 0 0.008f
r510 vdd_M2_3760_336 vdd_M2_3840_336 4.8
c1020 vdd_M2_3760_336 0 0.008f
c1021 vdd_M2_3840_336 0 0.008f
r511 vdd_M2_3840_336 vdd_M2_3920_336 4.8
c1022 vdd_M2_3840_336 0 0.008f
c1023 vdd_M2_3920_336 0 0.008f
r512 vdd_M2_3920_336 vdd_M2_3956_336 2.1599999999999997
c1024 vdd_M2_3920_336 0 0.0036f
c1025 vdd_M2_3956_336 0 0.0036f
r513 id_M2_364_252 id_M2_444_252 4.8
c1026 id_M2_364_252 0 0.008f
c1027 id_M2_444_252 0 0.008f
r514 id_M2_444_252 id_M2_524_252 4.8
c1028 id_M2_444_252 0 0.008f
c1029 id_M2_524_252 0 0.008f
r515 id_M2_524_252 id_M2_604_252 4.8
c1030 id_M2_524_252 0 0.008f
c1031 id_M2_604_252 0 0.008f
r516 id_M2_604_252 id_M2_684_252 4.8
c1032 id_M2_604_252 0 0.008f
c1033 id_M2_684_252 0 0.008f
r517 id_M2_684_252 id_M2_764_252 4.8
c1034 id_M2_684_252 0 0.008f
c1035 id_M2_764_252 0 0.008f
r518 id_M2_764_252 id_M2_844_252 4.8
c1036 id_M2_764_252 0 0.008f
c1037 id_M2_844_252 0 0.008f
r519 id_M2_844_252 id_M2_924_252 4.8
c1038 id_M2_844_252 0 0.008f
c1039 id_M2_924_252 0 0.008f
r520 id_M2_924_252 id_M2_1004_252 4.8
c1040 id_M2_924_252 0 0.008f
c1041 id_M2_1004_252 0 0.008f
r521 id_M2_1004_252 id_M2_1084_252 4.8
c1042 id_M2_1004_252 0 0.008f
c1043 id_M2_1084_252 0 0.008f
r522 id_M2_1084_252 id_M2_1164_252 4.8
c1044 id_M2_1084_252 0 0.008f
c1045 id_M2_1164_252 0 0.008f
r523 id_M2_1164_252 id_M2_1244_252 4.8
c1046 id_M2_1164_252 0 0.008f
c1047 id_M2_1244_252 0 0.008f
r524 id_M2_1244_252 id_M2_1324_252 4.8
c1048 id_M2_1244_252 0 0.008f
c1049 id_M2_1324_252 0 0.008f
r525 id_M2_1324_252 id_M2_1404_252 4.8
c1050 id_M2_1324_252 0 0.008f
c1051 id_M2_1404_252 0 0.008f
r526 id_M2_1404_252 id_M2_1484_252 4.8
c1052 id_M2_1404_252 0 0.008f
c1053 id_M2_1484_252 0 0.008f
r527 id_M2_1484_252 id_M2_1564_252 4.8
c1054 id_M2_1484_252 0 0.008f
c1055 id_M2_1564_252 0 0.008f
r528 id_M2_1564_252 id_M2_1644_252 4.8
c1056 id_M2_1564_252 0 0.008f
c1057 id_M2_1644_252 0 0.008f
r529 id_M2_1644_252 id_M2_1724_252 4.8
c1058 id_M2_1644_252 0 0.008f
c1059 id_M2_1724_252 0 0.008f
r530 id_M2_1724_252 id_M2_1804_252 4.8
c1060 id_M2_1724_252 0 0.008f
c1061 id_M2_1804_252 0 0.008f
r531 id_M2_1804_252 id_M2_1884_252 4.8
c1062 id_M2_1804_252 0 0.008f
c1063 id_M2_1884_252 0 0.008f
r532 id_M2_1884_252 id_M2_1964_252 4.8
c1064 id_M2_1884_252 0 0.008f
c1065 id_M2_1964_252 0 0.008f
r533 id_M2_1964_252 id_M2_2044_252 4.8
c1066 id_M2_1964_252 0 0.008f
c1067 id_M2_2044_252 0 0.008f
r534 id_M2_2044_252 id_M2_2124_252 4.8
c1068 id_M2_2044_252 0 0.008f
c1069 id_M2_2124_252 0 0.008f
r535 id_M2_2124_252 id_M2_2204_252 4.8
c1070 id_M2_2124_252 0 0.008f
c1071 id_M2_2204_252 0 0.008f
r536 id_M2_2204_252 id_M2_2284_252 4.8
c1072 id_M2_2204_252 0 0.008f
c1073 id_M2_2284_252 0 0.008f
r537 id_M2_2284_252 id_M2_2364_252 4.8
c1074 id_M2_2284_252 0 0.008f
c1075 id_M2_2364_252 0 0.008f
r538 id_M2_2364_252 id_M2_2444_252 4.8
c1076 id_M2_2364_252 0 0.008f
c1077 id_M2_2444_252 0 0.008f
r539 id_M2_2444_252 id_M2_2524_252 4.8
c1078 id_M2_2444_252 0 0.008f
c1079 id_M2_2524_252 0 0.008f
r540 id_M2_2524_252 id_M2_2604_252 4.8
c1080 id_M2_2524_252 0 0.008f
c1081 id_M2_2604_252 0 0.008f
r541 id_M2_2604_252 id_M2_2684_252 4.8
c1082 id_M2_2604_252 0 0.008f
c1083 id_M2_2684_252 0 0.008f
r542 id_M2_2684_252 id_M2_2764_252 4.8
c1084 id_M2_2684_252 0 0.008f
c1085 id_M2_2764_252 0 0.008f
r543 id_M2_2764_252 id_M2_2844_252 4.8
c1086 id_M2_2764_252 0 0.008f
c1087 id_M2_2844_252 0 0.008f
r544 id_M2_2844_252 id_M2_2924_252 4.8
c1088 id_M2_2844_252 0 0.008f
c1089 id_M2_2924_252 0 0.008f
r545 id_M2_2924_252 id_M2_3004_252 4.8
c1090 id_M2_2924_252 0 0.008f
c1091 id_M2_3004_252 0 0.008f
r546 id_M2_3004_252 id_M2_3084_252 4.8
c1092 id_M2_3004_252 0 0.008f
c1093 id_M2_3084_252 0 0.008f
r547 id_M2_3084_252 id_M2_3164_252 4.8
c1094 id_M2_3084_252 0 0.008f
c1095 id_M2_3164_252 0 0.008f
r548 id_M2_3164_252 id_M2_3244_252 4.8
c1096 id_M2_3164_252 0 0.008f
c1097 id_M2_3244_252 0 0.008f
r549 id_M2_3244_252 id_M2_3324_252 4.8
c1098 id_M2_3244_252 0 0.008f
c1099 id_M2_3324_252 0 0.008f
r550 id_M2_3324_252 id_M2_3404_252 4.8
c1100 id_M2_3324_252 0 0.008f
c1101 id_M2_3404_252 0 0.008f
r551 id_M2_3404_252 id_M2_3484_252 4.8
c1102 id_M2_3404_252 0 0.008f
c1103 id_M2_3484_252 0 0.008f
r552 id_M2_3484_252 id_M2_3564_252 4.8
c1104 id_M2_3484_252 0 0.008f
c1105 id_M2_3564_252 0 0.008f
r553 id_M2_3564_252 id_M2_3644_252 4.8
c1106 id_M2_3564_252 0 0.008f
c1107 id_M2_3644_252 0 0.008f
r554 id_M2_3644_252 id_M2_3724_252 4.8
c1108 id_M2_3644_252 0 0.008f
c1109 id_M2_3724_252 0 0.008f
r555 id_M2_3724_252 id_M2_3804_252 4.8
c1110 id_M2_3724_252 0 0.008f
c1111 id_M2_3804_252 0 0.008f
r556 id_M2_3804_252 id_M2_3840_252 2.1599999999999997
c1112 id_M2_3804_252 0 0.0036f
c1113 id_M2_3840_252 0 0.0036f
r557 vinp_M2_1324_252 vinp_M2_1404_252 4.8
c1114 vinp_M2_1324_252 0 0.008f
c1115 vinp_M2_1404_252 0 0.008f
r558 vinp_M2_1404_252 vinp_M2_1484_252 4.8
c1116 vinp_M2_1404_252 0 0.008f
c1117 vinp_M2_1484_252 0 0.008f
r559 vinp_M2_1484_252 vinp_M2_1564_252 4.8
c1118 vinp_M2_1484_252 0 0.008f
c1119 vinp_M2_1564_252 0 0.008f
r560 vinp_M2_1564_252 vinp_M2_1644_252 4.8
c1120 vinp_M2_1564_252 0 0.008f
c1121 vinp_M2_1644_252 0 0.008f
r561 vinp_M2_1644_252 vinp_M2_1724_252 4.8
c1122 vinp_M2_1644_252 0 0.008f
c1123 vinp_M2_1724_252 0 0.008f
r562 vinp_M2_1724_252 vinp_M2_1804_252 4.8
c1124 vinp_M2_1724_252 0 0.008f
c1125 vinp_M2_1804_252 0 0.008f
r563 vinp_M2_1804_252 vinp_M2_1884_252 4.8
c1126 vinp_M2_1804_252 0 0.008f
c1127 vinp_M2_1884_252 0 0.008f
r564 vinp_M2_1884_252 vinp_M2_1964_252 4.8
c1128 vinp_M2_1884_252 0 0.008f
c1129 vinp_M2_1964_252 0 0.008f
r565 vinp_M2_1964_252 vinp_M2_2044_252 4.8
c1130 vinp_M2_1964_252 0 0.008f
c1131 vinp_M2_2044_252 0 0.008f
r566 vinp_M2_2044_252 vinp_M2_2124_252 4.8
c1132 vinp_M2_2044_252 0 0.008f
c1133 vinp_M2_2124_252 0 0.008f
r567 vinp_M2_2124_252 vinp_M2_2204_252 4.8
c1134 vinp_M2_2124_252 0 0.008f
c1135 vinp_M2_2204_252 0 0.008f
r568 vinp_M2_2204_252 vinp_M2_2284_252 4.8
c1136 vinp_M2_2204_252 0 0.008f
c1137 vinp_M2_2284_252 0 0.008f
r569 vinp_M2_2284_252 vinp_M2_2364_252 4.8
c1138 vinp_M2_2284_252 0 0.008f
c1139 vinp_M2_2364_252 0 0.008f
r570 vinp_M2_2364_252 vinp_M2_2444_252 4.8
c1140 vinp_M2_2364_252 0 0.008f
c1141 vinp_M2_2444_252 0 0.008f
r571 vinp_M2_2444_252 vinp_M2_2524_252 4.8
c1142 vinp_M2_2444_252 0 0.008f
c1143 vinp_M2_2524_252 0 0.008f
r572 vinp_M2_2524_252 vinp_M2_2604_252 4.8
c1144 vinp_M2_2524_252 0 0.008f
c1145 vinp_M2_2604_252 0 0.008f
r573 vinp_M2_2604_252 vinp_M2_2684_252 4.8
c1146 vinp_M2_2604_252 0 0.008f
c1147 vinp_M2_2684_252 0 0.008f
r574 vinp_M2_2684_252 vinp_M2_2764_252 4.8
c1148 vinp_M2_2684_252 0 0.008f
c1149 vinp_M2_2764_252 0 0.008f
r575 vinp_M2_2764_252 vinp_M2_2844_252 4.8
c1150 vinp_M2_2764_252 0 0.008f
c1151 vinp_M2_2844_252 0 0.008f
r576 vinp_M2_2844_252 vinp_M2_2924_252 4.8
c1152 vinp_M2_2844_252 0 0.008f
c1153 vinp_M2_2924_252 0 0.008f
r577 vinp_M2_2924_252 vinp_M2_3004_252 4.8
c1154 vinp_M2_2924_252 0 0.008f
c1155 vinp_M2_3004_252 0 0.008f
r578 vinp_M2_3004_252 vinp_M2_3084_252 4.8
c1156 vinp_M2_3004_252 0 0.008f
c1157 vinp_M2_3084_252 0 0.008f
r579 vinp_M2_3084_252 vinp_M2_3164_252 4.8
c1158 vinp_M2_3084_252 0 0.008f
c1159 vinp_M2_3164_252 0 0.008f
r580 vinp_M2_3164_252 vinp_M2_3244_252 4.8
c1160 vinp_M2_3164_252 0 0.008f
c1161 vinp_M2_3244_252 0 0.008f
r581 vinp_M2_3244_252 vinp_M2_3324_252 4.8
c1162 vinp_M2_3244_252 0 0.008f
c1163 vinp_M2_3324_252 0 0.008f
r582 vinp_M2_3324_252 vinp_M2_3404_252 4.8
c1164 vinp_M2_3324_252 0 0.008f
c1165 vinp_M2_3404_252 0 0.008f
r583 vinp_M2_3404_252 vinp_M2_3484_252 4.8
c1166 vinp_M2_3404_252 0 0.008f
c1167 vinp_M2_3484_252 0 0.008f
r584 vinp_M2_3484_252 vinp_M2_3564_252 4.8
c1168 vinp_M2_3484_252 0 0.008f
c1169 vinp_M2_3564_252 0 0.008f
r585 vinp_M2_3564_252 vinp_M2_3644_252 4.8
c1170 vinp_M2_3564_252 0 0.008f
c1171 vinp_M2_3644_252 0 0.008f
r586 vinp_M2_3644_252 vinp_M2_3724_252 4.8
c1172 vinp_M2_3644_252 0 0.008f
c1173 vinp_M2_3724_252 0 0.008f
r587 vinp_M2_3724_252 vinp_M2_3804_252 4.8
c1174 vinp_M2_3724_252 0 0.008f
c1175 vinp_M2_3804_252 0 0.008f
r588 vinp_M2_3804_252 vinp_M2_3840_252 2.1599999999999997
c1176 vinp_M2_3804_252 0 0.0036f
c1177 vinp_M2_3840_252 0 0.0036f
r589 net8_M2_1804_252 net8_M2_1884_252 4.8
c1178 net8_M2_1804_252 0 0.008f
c1179 net8_M2_1884_252 0 0.008f
r590 net8_M2_1884_252 net8_M2_1964_252 4.8
c1180 net8_M2_1884_252 0 0.008f
c1181 net8_M2_1964_252 0 0.008f
r591 net8_M2_1964_252 net8_M2_2044_252 4.8
c1182 net8_M2_1964_252 0 0.008f
c1183 net8_M2_2044_252 0 0.008f
r592 net8_M2_2044_252 net8_M2_2124_252 4.8
c1184 net8_M2_2044_252 0 0.008f
c1185 net8_M2_2124_252 0 0.008f
r593 net8_M2_2124_252 net8_M2_2204_252 4.8
c1186 net8_M2_2124_252 0 0.008f
c1187 net8_M2_2204_252 0 0.008f
r594 net8_M2_2204_252 net8_M2_2284_252 4.8
c1188 net8_M2_2204_252 0 0.008f
c1189 net8_M2_2284_252 0 0.008f
r595 net8_M2_2284_252 net8_M2_2364_252 4.8
c1190 net8_M2_2284_252 0 0.008f
c1191 net8_M2_2364_252 0 0.008f
r596 net8_M2_2364_252 net8_M2_2444_252 4.8
c1192 net8_M2_2364_252 0 0.008f
c1193 net8_M2_2444_252 0 0.008f
r597 net8_M2_2444_252 net8_M2_2524_252 4.8
c1194 net8_M2_2444_252 0 0.008f
c1195 net8_M2_2524_252 0 0.008f
r598 net8_M2_2524_252 net8_M2_2604_252 4.8
c1196 net8_M2_2524_252 0 0.008f
c1197 net8_M2_2604_252 0 0.008f
r599 net8_M2_2604_252 net8_M2_2684_252 4.8
c1198 net8_M2_2604_252 0 0.008f
c1199 net8_M2_2684_252 0 0.008f
r600 net8_M2_2684_252 net8_M2_2764_252 4.8
c1200 net8_M2_2684_252 0 0.008f
c1201 net8_M2_2764_252 0 0.008f
r601 net8_M2_2764_252 net8_M2_2844_252 4.8
c1202 net8_M2_2764_252 0 0.008f
c1203 net8_M2_2844_252 0 0.008f
r602 net8_M2_2844_252 net8_M2_2924_252 4.8
c1204 net8_M2_2844_252 0 0.008f
c1205 net8_M2_2924_252 0 0.008f
r603 net8_M2_2924_252 net8_M2_3004_252 4.8
c1206 net8_M2_2924_252 0 0.008f
c1207 net8_M2_3004_252 0 0.008f
r604 net8_M2_3004_252 net8_M2_3084_252 4.8
c1208 net8_M2_3004_252 0 0.008f
c1209 net8_M2_3084_252 0 0.008f
r605 net8_M2_3084_252 net8_M2_3164_252 4.8
c1210 net8_M2_3084_252 0 0.008f
c1211 net8_M2_3164_252 0 0.008f
r606 net8_M2_3164_252 net8_M2_3244_252 4.8
c1212 net8_M2_3164_252 0 0.008f
c1213 net8_M2_3244_252 0 0.008f
r607 net8_M2_3244_252 net8_M2_3324_252 4.8
c1214 net8_M2_3244_252 0 0.008f
c1215 net8_M2_3324_252 0 0.008f
r608 net8_M2_3324_252 net8_M2_3404_252 4.8
c1216 net8_M2_3324_252 0 0.008f
c1217 net8_M2_3404_252 0 0.008f
r609 net8_M2_3404_252 net8_M2_3484_252 4.8
c1218 net8_M2_3404_252 0 0.008f
c1219 net8_M2_3484_252 0 0.008f
r610 net8_M2_3484_252 net8_M2_3564_252 4.8
c1220 net8_M2_3484_252 0 0.008f
c1221 net8_M2_3564_252 0 0.008f
r611 net8_M2_3564_252 net8_M2_3644_252 4.8
c1222 net8_M2_3564_252 0 0.008f
c1223 net8_M2_3644_252 0 0.008f
r612 net8_M2_3644_252 net8_M2_3724_252 4.8
c1224 net8_M2_3644_252 0 0.008f
c1225 net8_M2_3724_252 0 0.008f
r613 net8_M2_3724_252 net8_M2_3804_252 4.8
c1226 net8_M2_3724_252 0 0.008f
c1227 net8_M2_3804_252 0 0.008f
r614 net8_M2_3804_252 net8_M2_3840_252 2.1599999999999997
c1228 net8_M2_3804_252 0 0.0036f
c1229 net8_M2_3840_252 0 0.0036f
r615 vout_M2_2364_252 vout_M2_2444_252 4.8
c1230 vout_M2_2364_252 0 0.008f
c1231 vout_M2_2444_252 0 0.008f
r616 vout_M2_2444_252 vout_M2_2524_252 4.8
c1232 vout_M2_2444_252 0 0.008f
c1233 vout_M2_2524_252 0 0.008f
r617 vout_M2_2524_252 vout_M2_2604_252 4.8
c1234 vout_M2_2524_252 0 0.008f
c1235 vout_M2_2604_252 0 0.008f
r618 vout_M2_2604_252 vout_M2_2684_252 4.8
c1236 vout_M2_2604_252 0 0.008f
c1237 vout_M2_2684_252 0 0.008f
r619 vout_M2_2684_252 vout_M2_2764_252 4.8
c1238 vout_M2_2684_252 0 0.008f
c1239 vout_M2_2764_252 0 0.008f
r620 vout_M2_2764_252 vout_M2_2844_252 4.8
c1240 vout_M2_2764_252 0 0.008f
c1241 vout_M2_2844_252 0 0.008f
r621 vout_M2_2844_252 vout_M2_2924_252 4.8
c1242 vout_M2_2844_252 0 0.008f
c1243 vout_M2_2924_252 0 0.008f
r622 vout_M2_2924_252 vout_M2_3004_252 4.8
c1244 vout_M2_2924_252 0 0.008f
c1245 vout_M2_3004_252 0 0.008f
r623 vout_M2_3004_252 vout_M2_3084_252 4.8
c1246 vout_M2_3004_252 0 0.008f
c1247 vout_M2_3084_252 0 0.008f
r624 vout_M2_3084_252 vout_M2_3164_252 4.8
c1248 vout_M2_3084_252 0 0.008f
c1249 vout_M2_3164_252 0 0.008f
r625 vout_M2_3164_252 vout_M2_3244_252 4.8
c1250 vout_M2_3164_252 0 0.008f
c1251 vout_M2_3244_252 0 0.008f
r626 vout_M2_3244_252 vout_M2_3324_252 4.8
c1252 vout_M2_3244_252 0 0.008f
c1253 vout_M2_3324_252 0 0.008f
r627 vout_M2_3324_252 vout_M2_3404_252 4.8
c1254 vout_M2_3324_252 0 0.008f
c1255 vout_M2_3404_252 0 0.008f
r628 vout_M2_3404_252 vout_M2_3484_252 4.8
c1256 vout_M2_3404_252 0 0.008f
c1257 vout_M2_3484_252 0 0.008f
r629 vout_M2_3484_252 vout_M2_3564_252 4.8
c1258 vout_M2_3484_252 0 0.008f
c1259 vout_M2_3564_252 0 0.008f
r630 vout_M2_3564_252 vout_M2_3644_252 4.8
c1260 vout_M2_3564_252 0 0.008f
c1261 vout_M2_3644_252 0 0.008f
r631 vout_M2_3644_252 vout_M2_3724_252 4.8
c1262 vout_M2_3644_252 0 0.008f
c1263 vout_M2_3724_252 0 0.008f
r632 vout_M2_3724_252 vout_M2_3804_252 4.8
c1264 vout_M2_3724_252 0 0.008f
c1265 vout_M2_3804_252 0 0.008f
r633 vout_M2_3804_252 vout_M2_3840_252 2.1599999999999997
c1266 vout_M2_3804_252 0 0.0036f
c1267 vout_M2_3840_252 0 0.0036f
r634 net8_M2_400_252 net8_M2_480_252 4.8
c1268 net8_M2_400_252 0 0.008f
c1269 net8_M2_480_252 0 0.008f
r635 net8_M2_480_252 net8_M2_560_252 4.8
c1270 net8_M2_480_252 0 0.008f
c1271 net8_M2_560_252 0 0.008f
r636 net8_M2_560_252 net8_M2_640_252 4.8
c1272 net8_M2_560_252 0 0.008f
c1273 net8_M2_640_252 0 0.008f
r637 net8_M2_640_252 net8_M2_720_252 4.8
c1274 net8_M2_640_252 0 0.008f
c1275 net8_M2_720_252 0 0.008f
r638 net8_M2_720_252 net8_M2_800_252 4.8
c1276 net8_M2_720_252 0 0.008f
c1277 net8_M2_800_252 0 0.008f
r639 net8_M2_800_252 net8_M2_880_252 4.8
c1278 net8_M2_800_252 0 0.008f
c1279 net8_M2_880_252 0 0.008f
r640 net8_M2_880_252 net8_M2_960_252 4.8
c1280 net8_M2_880_252 0 0.008f
c1281 net8_M2_960_252 0 0.008f
r641 net8_M2_960_252 net8_M2_1040_252 4.8
c1282 net8_M2_960_252 0 0.008f
c1283 net8_M2_1040_252 0 0.008f
r642 net8_M2_1040_252 net8_M2_1120_252 4.8
c1284 net8_M2_1040_252 0 0.008f
c1285 net8_M2_1120_252 0 0.008f
r643 net8_M2_1120_252 net8_M2_1200_252 4.8
c1286 net8_M2_1120_252 0 0.008f
c1287 net8_M2_1200_252 0 0.008f
r644 net8_M2_1200_252 net8_M2_1280_252 4.8
c1288 net8_M2_1200_252 0 0.008f
c1289 net8_M2_1280_252 0 0.008f
r645 net8_M2_1280_252 net8_M2_1360_252 4.8
c1290 net8_M2_1280_252 0 0.008f
c1291 net8_M2_1360_252 0 0.008f
r646 net8_M2_1360_252 net8_M2_1440_252 4.8
c1292 net8_M2_1360_252 0 0.008f
c1293 net8_M2_1440_252 0 0.008f
r647 net8_M2_1440_252 net8_M2_1520_252 4.8
c1294 net8_M2_1440_252 0 0.008f
c1295 net8_M2_1520_252 0 0.008f
r648 net8_M2_1520_252 net8_M2_1600_252 4.8
c1296 net8_M2_1520_252 0 0.008f
c1297 net8_M2_1600_252 0 0.008f
r649 net8_M2_1600_252 net8_M2_1680_252 4.8
c1298 net8_M2_1600_252 0 0.008f
c1299 net8_M2_1680_252 0 0.008f
r650 net8_M2_1680_252 net8_M2_1760_252 4.8
c1300 net8_M2_1680_252 0 0.008f
c1301 net8_M2_1760_252 0 0.008f
r651 net8_M2_1760_252 net8_M2_1840_252 4.8
c1302 net8_M2_1760_252 0 0.008f
c1303 net8_M2_1840_252 0 0.008f
r652 net8_M2_1840_252 net8_M2_1920_252 4.8
c1304 net8_M2_1840_252 0 0.008f
c1305 net8_M2_1920_252 0 0.008f
r653 net8_M2_1920_252 net8_M2_2000_252 4.8
c1306 net8_M2_1920_252 0 0.008f
c1307 net8_M2_2000_252 0 0.008f
r654 net8_M2_2000_252 net8_M2_2080_252 4.8
c1308 net8_M2_2000_252 0 0.008f
c1309 net8_M2_2080_252 0 0.008f
r655 net8_M2_2080_252 net8_M2_2160_252 4.8
c1310 net8_M2_2080_252 0 0.008f
c1311 net8_M2_2160_252 0 0.008f
r656 net8_M2_2160_252 net8_M2_2240_252 4.8
c1312 net8_M2_2160_252 0 0.008f
c1313 net8_M2_2240_252 0 0.008f
r657 net8_M2_2240_252 net8_M2_2320_252 4.8
c1314 net8_M2_2240_252 0 0.008f
c1315 net8_M2_2320_252 0 0.008f
r658 net8_M2_2320_252 net8_M2_2400_252 4.8
c1316 net8_M2_2320_252 0 0.008f
c1317 net8_M2_2400_252 0 0.008f
r659 net8_M2_2400_252 net8_M2_2480_252 4.8
c1318 net8_M2_2400_252 0 0.008f
c1319 net8_M2_2480_252 0 0.008f
r660 net8_M2_2480_252 net8_M2_2560_252 4.8
c1320 net8_M2_2480_252 0 0.008f
c1321 net8_M2_2560_252 0 0.008f
r661 net8_M2_2560_252 net8_M2_2640_252 4.8
c1322 net8_M2_2560_252 0 0.008f
c1323 net8_M2_2640_252 0 0.008f
r662 net8_M2_2640_252 net8_M2_2720_252 4.8
c1324 net8_M2_2640_252 0 0.008f
c1325 net8_M2_2720_252 0 0.008f
r663 net8_M2_2720_252 net8_M2_2800_252 4.8
c1326 net8_M2_2720_252 0 0.008f
c1327 net8_M2_2800_252 0 0.008f
r664 net8_M2_2800_252 net8_M2_2880_252 4.8
c1328 net8_M2_2800_252 0 0.008f
c1329 net8_M2_2880_252 0 0.008f
r665 net8_M2_2880_252 net8_M2_2960_252 4.8
c1330 net8_M2_2880_252 0 0.008f
c1331 net8_M2_2960_252 0 0.008f
r666 net8_M2_2960_252 net8_M2_3040_252 4.8
c1332 net8_M2_2960_252 0 0.008f
c1333 net8_M2_3040_252 0 0.008f
r667 net8_M2_3040_252 net8_M2_3120_252 4.8
c1334 net8_M2_3040_252 0 0.008f
c1335 net8_M2_3120_252 0 0.008f
r668 net8_M2_3120_252 net8_M2_3200_252 4.8
c1336 net8_M2_3120_252 0 0.008f
c1337 net8_M2_3200_252 0 0.008f
r669 net8_M2_3200_252 net8_M2_3280_252 4.8
c1338 net8_M2_3200_252 0 0.008f
c1339 net8_M2_3280_252 0 0.008f
r670 net8_M2_3280_252 net8_M2_3360_252 4.8
c1340 net8_M2_3280_252 0 0.008f
c1341 net8_M2_3360_252 0 0.008f
r671 net8_M2_3360_252 net8_M2_3440_252 4.8
c1342 net8_M2_3360_252 0 0.008f
c1343 net8_M2_3440_252 0 0.008f
r672 net8_M2_3440_252 net8_M2_3520_252 4.8
c1344 net8_M2_3440_252 0 0.008f
c1345 net8_M2_3520_252 0 0.008f
r673 net8_M2_3520_252 net8_M2_3600_252 4.8
c1346 net8_M2_3520_252 0 0.008f
c1347 net8_M2_3600_252 0 0.008f
r674 net8_M2_3600_252 net8_M2_3680_252 4.8
c1348 net8_M2_3600_252 0 0.008f
c1349 net8_M2_3680_252 0 0.008f
r675 net8_M2_3680_252 net8_M2_3760_252 4.8
c1350 net8_M2_3680_252 0 0.008f
c1351 net8_M2_3760_252 0 0.008f
r676 net8_M2_3760_252 net8_M2_3840_252 4.8
c1352 net8_M2_3760_252 0 0.008f
c1353 net8_M2_3840_252 0 0.008f
r677 net8_M2_3840_252 net8_M2_3920_252 4.8
c1354 net8_M2_3840_252 0 0.008f
c1355 net8_M2_3920_252 0 0.008f
r678 net8_M2_3920_252 net8_M2_3956_252 2.1599999999999997
c1356 net8_M2_3920_252 0 0.0036f
c1357 net8_M2_3956_252 0 0.0036f
r679 vss_M2_284_420 vss_M2_364_420 4.8
c1358 vss_M2_284_420 0 0.008f
c1359 vss_M2_364_420 0 0.008f
r680 vss_M2_364_420 vss_M2_444_420 4.8
c1360 vss_M2_364_420 0 0.008f
c1361 vss_M2_444_420 0 0.008f
r681 vss_M2_444_420 vss_M2_524_420 4.8
c1362 vss_M2_444_420 0 0.008f
c1363 vss_M2_524_420 0 0.008f
r682 vss_M2_524_420 vss_M2_604_420 4.8
c1364 vss_M2_524_420 0 0.008f
c1365 vss_M2_604_420 0 0.008f
r683 vss_M2_604_420 vss_M2_684_420 4.8
c1366 vss_M2_604_420 0 0.008f
c1367 vss_M2_684_420 0 0.008f
r684 vss_M2_684_420 vss_M2_764_420 4.8
c1368 vss_M2_684_420 0 0.008f
c1369 vss_M2_764_420 0 0.008f
r685 vss_M2_764_420 vss_M2_844_420 4.8
c1370 vss_M2_764_420 0 0.008f
c1371 vss_M2_844_420 0 0.008f
r686 vss_M2_844_420 vss_M2_924_420 4.8
c1372 vss_M2_844_420 0 0.008f
c1373 vss_M2_924_420 0 0.008f
r687 vss_M2_924_420 vss_M2_1004_420 4.8
c1374 vss_M2_924_420 0 0.008f
c1375 vss_M2_1004_420 0 0.008f
r688 vss_M2_1004_420 vss_M2_1084_420 4.8
c1376 vss_M2_1004_420 0 0.008f
c1377 vss_M2_1084_420 0 0.008f
r689 vss_M2_1084_420 vss_M2_1164_420 4.8
c1378 vss_M2_1084_420 0 0.008f
c1379 vss_M2_1164_420 0 0.008f
r690 vss_M2_1164_420 vss_M2_1244_420 4.8
c1380 vss_M2_1164_420 0 0.008f
c1381 vss_M2_1244_420 0 0.008f
r691 vss_M2_1244_420 vss_M2_1324_420 4.8
c1382 vss_M2_1244_420 0 0.008f
c1383 vss_M2_1324_420 0 0.008f
r692 vss_M2_1324_420 vss_M2_1404_420 4.8
c1384 vss_M2_1324_420 0 0.008f
c1385 vss_M2_1404_420 0 0.008f
r693 vss_M2_1404_420 vss_M2_1484_420 4.8
c1386 vss_M2_1404_420 0 0.008f
c1387 vss_M2_1484_420 0 0.008f
r694 vss_M2_1484_420 vss_M2_1564_420 4.8
c1388 vss_M2_1484_420 0 0.008f
c1389 vss_M2_1564_420 0 0.008f
r695 vss_M2_1564_420 vss_M2_1644_420 4.8
c1390 vss_M2_1564_420 0 0.008f
c1391 vss_M2_1644_420 0 0.008f
r696 vss_M2_1644_420 vss_M2_1724_420 4.8
c1392 vss_M2_1644_420 0 0.008f
c1393 vss_M2_1724_420 0 0.008f
r697 vss_M2_1724_420 vss_M2_1804_420 4.8
c1394 vss_M2_1724_420 0 0.008f
c1395 vss_M2_1804_420 0 0.008f
r698 vss_M2_1804_420 vss_M2_1884_420 4.8
c1396 vss_M2_1804_420 0 0.008f
c1397 vss_M2_1884_420 0 0.008f
r699 vss_M2_1884_420 vss_M2_1964_420 4.8
c1398 vss_M2_1884_420 0 0.008f
c1399 vss_M2_1964_420 0 0.008f
r700 vss_M2_1964_420 vss_M2_2044_420 4.8
c1400 vss_M2_1964_420 0 0.008f
c1401 vss_M2_2044_420 0 0.008f
r701 vss_M2_2044_420 vss_M2_2124_420 4.8
c1402 vss_M2_2044_420 0 0.008f
c1403 vss_M2_2124_420 0 0.008f
r702 vss_M2_2124_420 vss_M2_2204_420 4.8
c1404 vss_M2_2124_420 0 0.008f
c1405 vss_M2_2204_420 0 0.008f
r703 vss_M2_2204_420 vss_M2_2284_420 4.8
c1406 vss_M2_2204_420 0 0.008f
c1407 vss_M2_2284_420 0 0.008f
r704 vss_M2_2284_420 vss_M2_2364_420 4.8
c1408 vss_M2_2284_420 0 0.008f
c1409 vss_M2_2364_420 0 0.008f
r705 vss_M2_2364_420 vss_M2_2444_420 4.8
c1410 vss_M2_2364_420 0 0.008f
c1411 vss_M2_2444_420 0 0.008f
r706 vss_M2_2444_420 vss_M2_2524_420 4.8
c1412 vss_M2_2444_420 0 0.008f
c1413 vss_M2_2524_420 0 0.008f
r707 vss_M2_2524_420 vss_M2_2604_420 4.8
c1414 vss_M2_2524_420 0 0.008f
c1415 vss_M2_2604_420 0 0.008f
r708 vss_M2_2604_420 vss_M2_2684_420 4.8
c1416 vss_M2_2604_420 0 0.008f
c1417 vss_M2_2684_420 0 0.008f
r709 vss_M2_2684_420 vss_M2_2764_420 4.8
c1418 vss_M2_2684_420 0 0.008f
c1419 vss_M2_2764_420 0 0.008f
r710 vss_M2_2764_420 vss_M2_2844_420 4.8
c1420 vss_M2_2764_420 0 0.008f
c1421 vss_M2_2844_420 0 0.008f
r711 vss_M2_2844_420 vss_M2_2924_420 4.8
c1422 vss_M2_2844_420 0 0.008f
c1423 vss_M2_2924_420 0 0.008f
r712 vss_M2_2924_420 vss_M2_3004_420 4.8
c1424 vss_M2_2924_420 0 0.008f
c1425 vss_M2_3004_420 0 0.008f
r713 vss_M2_3004_420 vss_M2_3084_420 4.8
c1426 vss_M2_3004_420 0 0.008f
c1427 vss_M2_3084_420 0 0.008f
r714 vss_M2_3084_420 vss_M2_3164_420 4.8
c1428 vss_M2_3084_420 0 0.008f
c1429 vss_M2_3164_420 0 0.008f
r715 vss_M2_3164_420 vss_M2_3244_420 4.8
c1430 vss_M2_3164_420 0 0.008f
c1431 vss_M2_3244_420 0 0.008f
r716 vss_M2_3244_420 vss_M2_3324_420 4.8
c1432 vss_M2_3244_420 0 0.008f
c1433 vss_M2_3324_420 0 0.008f
r717 vss_M2_3324_420 vss_M2_3404_420 4.8
c1434 vss_M2_3324_420 0 0.008f
c1435 vss_M2_3404_420 0 0.008f
r718 vss_M2_3404_420 vss_M2_3484_420 4.8
c1436 vss_M2_3404_420 0 0.008f
c1437 vss_M2_3484_420 0 0.008f
r719 vss_M2_3484_420 vss_M2_3564_420 4.8
c1438 vss_M2_3484_420 0 0.008f
c1439 vss_M2_3564_420 0 0.008f
r720 vss_M2_3564_420 vss_M2_3644_420 4.8
c1440 vss_M2_3564_420 0 0.008f
c1441 vss_M2_3644_420 0 0.008f
r721 vss_M2_3644_420 vss_M2_3724_420 4.8
c1442 vss_M2_3644_420 0 0.008f
c1443 vss_M2_3724_420 0 0.008f
r722 vss_M2_3724_420 vss_M2_3804_420 4.8
c1444 vss_M2_3724_420 0 0.008f
c1445 vss_M2_3804_420 0 0.008f
r723 vss_M2_3804_420 vss_M2_3840_420 2.1599999999999997
c1446 vss_M2_3804_420 0 0.0036f
c1447 vss_M2_3840_420 0 0.0036f
r724 vinp_M2_1724_420 vinp_M2_1804_420 4.8
c1448 vinp_M2_1724_420 0 0.008f
c1449 vinp_M2_1804_420 0 0.008f
r725 vinp_M2_1804_420 vinp_M2_1884_420 4.8
c1450 vinp_M2_1804_420 0 0.008f
c1451 vinp_M2_1884_420 0 0.008f
r726 vinp_M2_1884_420 vinp_M2_1964_420 4.8
c1452 vinp_M2_1884_420 0 0.008f
c1453 vinp_M2_1964_420 0 0.008f
r727 vinp_M2_1964_420 vinp_M2_2044_420 4.8
c1454 vinp_M2_1964_420 0 0.008f
c1455 vinp_M2_2044_420 0 0.008f
r728 vinp_M2_2044_420 vinp_M2_2124_420 4.8
c1456 vinp_M2_2044_420 0 0.008f
c1457 vinp_M2_2124_420 0 0.008f
r729 vinp_M2_2124_420 vinp_M2_2204_420 4.8
c1458 vinp_M2_2124_420 0 0.008f
c1459 vinp_M2_2204_420 0 0.008f
r730 vinp_M2_2204_420 vinp_M2_2284_420 4.8
c1460 vinp_M2_2204_420 0 0.008f
c1461 vinp_M2_2284_420 0 0.008f
r731 vinp_M2_2284_420 vinp_M2_2364_420 4.8
c1462 vinp_M2_2284_420 0 0.008f
c1463 vinp_M2_2364_420 0 0.008f
r732 vinp_M2_2364_420 vinp_M2_2444_420 4.8
c1464 vinp_M2_2364_420 0 0.008f
c1465 vinp_M2_2444_420 0 0.008f
r733 vinp_M2_2444_420 vinp_M2_2524_420 4.8
c1466 vinp_M2_2444_420 0 0.008f
c1467 vinp_M2_2524_420 0 0.008f
r734 vinp_M2_2524_420 vinp_M2_2604_420 4.8
c1468 vinp_M2_2524_420 0 0.008f
c1469 vinp_M2_2604_420 0 0.008f
r735 vinp_M2_2604_420 vinp_M2_2684_420 4.8
c1470 vinp_M2_2604_420 0 0.008f
c1471 vinp_M2_2684_420 0 0.008f
r736 vinp_M2_2684_420 vinp_M2_2764_420 4.8
c1472 vinp_M2_2684_420 0 0.008f
c1473 vinp_M2_2764_420 0 0.008f
r737 vinp_M2_2764_420 vinp_M2_2844_420 4.8
c1474 vinp_M2_2764_420 0 0.008f
c1475 vinp_M2_2844_420 0 0.008f
r738 vinp_M2_2844_420 vinp_M2_2924_420 4.8
c1476 vinp_M2_2844_420 0 0.008f
c1477 vinp_M2_2924_420 0 0.008f
r739 vinp_M2_2924_420 vinp_M2_3004_420 4.8
c1478 vinp_M2_2924_420 0 0.008f
c1479 vinp_M2_3004_420 0 0.008f
r740 vinp_M2_3004_420 vinp_M2_3084_420 4.8
c1480 vinp_M2_3004_420 0 0.008f
c1481 vinp_M2_3084_420 0 0.008f
r741 vinp_M2_3084_420 vinp_M2_3164_420 4.8
c1482 vinp_M2_3084_420 0 0.008f
c1483 vinp_M2_3164_420 0 0.008f
r742 vinp_M2_3164_420 vinp_M2_3244_420 4.8
c1484 vinp_M2_3164_420 0 0.008f
c1485 vinp_M2_3244_420 0 0.008f
r743 vinp_M2_3244_420 vinp_M2_3324_420 4.8
c1486 vinp_M2_3244_420 0 0.008f
c1487 vinp_M2_3324_420 0 0.008f
r744 vinp_M2_3324_420 vinp_M2_3404_420 4.8
c1488 vinp_M2_3324_420 0 0.008f
c1489 vinp_M2_3404_420 0 0.008f
r745 vinp_M2_3404_420 vinp_M2_3484_420 4.8
c1490 vinp_M2_3404_420 0 0.008f
c1491 vinp_M2_3484_420 0 0.008f
r746 vinp_M2_3484_420 vinp_M2_3564_420 4.8
c1492 vinp_M2_3484_420 0 0.008f
c1493 vinp_M2_3564_420 0 0.008f
r747 vinp_M2_3564_420 vinp_M2_3644_420 4.8
c1494 vinp_M2_3564_420 0 0.008f
c1495 vinp_M2_3644_420 0 0.008f
r748 vinp_M2_3644_420 vinp_M2_3724_420 4.8
c1496 vinp_M2_3644_420 0 0.008f
c1497 vinp_M2_3724_420 0 0.008f
r749 vinp_M2_3724_420 vinp_M2_3804_420 4.8
c1498 vinp_M2_3724_420 0 0.008f
c1499 vinp_M2_3804_420 0 0.008f
r750 vinp_M2_3804_420 vinp_M2_3840_420 2.1599999999999997
c1500 vinp_M2_3804_420 0 0.0036f
c1501 vinp_M2_3840_420 0 0.0036f
r751 vdd_M2_3004_420 vdd_M2_3084_420 4.8
c1502 vdd_M2_3004_420 0 0.008f
c1503 vdd_M2_3084_420 0 0.008f
r752 vdd_M2_3084_420 vdd_M2_3164_420 4.8
c1504 vdd_M2_3084_420 0 0.008f
c1505 vdd_M2_3164_420 0 0.008f
r753 vdd_M2_3164_420 vdd_M2_3244_420 4.8
c1506 vdd_M2_3164_420 0 0.008f
c1507 vdd_M2_3244_420 0 0.008f
r754 vdd_M2_3244_420 vdd_M2_3324_420 4.8
c1508 vdd_M2_3244_420 0 0.008f
c1509 vdd_M2_3324_420 0 0.008f
r755 vdd_M2_3324_420 vdd_M2_3404_420 4.8
c1510 vdd_M2_3324_420 0 0.008f
c1511 vdd_M2_3404_420 0 0.008f
r756 vdd_M2_3404_420 vdd_M2_3484_420 4.8
c1512 vdd_M2_3404_420 0 0.008f
c1513 vdd_M2_3484_420 0 0.008f
r757 vdd_M2_3484_420 vdd_M2_3564_420 4.8
c1514 vdd_M2_3484_420 0 0.008f
c1515 vdd_M2_3564_420 0 0.008f
r758 vdd_M2_3564_420 vdd_M2_3644_420 4.8
c1516 vdd_M2_3564_420 0 0.008f
c1517 vdd_M2_3644_420 0 0.008f
r759 vdd_M2_3644_420 vdd_M2_3724_420 4.8
c1518 vdd_M2_3644_420 0 0.008f
c1519 vdd_M2_3724_420 0 0.008f
r760 vdd_M2_3724_420 vdd_M2_3804_420 4.8
c1520 vdd_M2_3724_420 0 0.008f
c1521 vdd_M2_3804_420 0 0.008f
r761 vdd_M2_3804_420 vdd_M2_3840_420 2.1599999999999997
c1522 vdd_M2_3804_420 0 0.0036f
c1523 vdd_M2_3840_420 0 0.0036f
r762 net8_M2_3644_420 net8_M2_3724_420 4.8
c1524 net8_M2_3644_420 0 0.008f
c1525 net8_M2_3724_420 0 0.008f
r763 net8_M2_3724_420 net8_M2_3804_420 4.8
c1526 net8_M2_3724_420 0 0.008f
c1527 net8_M2_3804_420 0 0.008f
r764 net8_M2_3804_420 net8_M2_3840_420 2.1599999999999997
c1528 net8_M2_3804_420 0 0.0036f
c1529 net8_M2_3840_420 0 0.0036f
r765 net8_M2_320_420 net8_M2_400_420 4.8
c1530 net8_M2_320_420 0 0.008f
c1531 net8_M2_400_420 0 0.008f
r766 net8_M2_400_420 net8_M2_480_420 4.8
c1532 net8_M2_400_420 0 0.008f
c1533 net8_M2_480_420 0 0.008f
r767 net8_M2_480_420 net8_M2_560_420 4.8
c1534 net8_M2_480_420 0 0.008f
c1535 net8_M2_560_420 0 0.008f
r768 net8_M2_560_420 net8_M2_640_420 4.8
c1536 net8_M2_560_420 0 0.008f
c1537 net8_M2_640_420 0 0.008f
r769 net8_M2_640_420 net8_M2_720_420 4.8
c1538 net8_M2_640_420 0 0.008f
c1539 net8_M2_720_420 0 0.008f
r770 net8_M2_720_420 net8_M2_800_420 4.8
c1540 net8_M2_720_420 0 0.008f
c1541 net8_M2_800_420 0 0.008f
r771 net8_M2_800_420 net8_M2_880_420 4.8
c1542 net8_M2_800_420 0 0.008f
c1543 net8_M2_880_420 0 0.008f
r772 net8_M2_880_420 net8_M2_960_420 4.8
c1544 net8_M2_880_420 0 0.008f
c1545 net8_M2_960_420 0 0.008f
r773 net8_M2_960_420 net8_M2_1040_420 4.8
c1546 net8_M2_960_420 0 0.008f
c1547 net8_M2_1040_420 0 0.008f
r774 net8_M2_1040_420 net8_M2_1120_420 4.8
c1548 net8_M2_1040_420 0 0.008f
c1549 net8_M2_1120_420 0 0.008f
r775 net8_M2_1120_420 net8_M2_1200_420 4.8
c1550 net8_M2_1120_420 0 0.008f
c1551 net8_M2_1200_420 0 0.008f
r776 net8_M2_1200_420 net8_M2_1280_420 4.8
c1552 net8_M2_1200_420 0 0.008f
c1553 net8_M2_1280_420 0 0.008f
r777 net8_M2_1280_420 net8_M2_1360_420 4.8
c1554 net8_M2_1280_420 0 0.008f
c1555 net8_M2_1360_420 0 0.008f
r778 net8_M2_1360_420 net8_M2_1440_420 4.8
c1556 net8_M2_1360_420 0 0.008f
c1557 net8_M2_1440_420 0 0.008f
r779 net8_M2_1440_420 net8_M2_1520_420 4.8
c1558 net8_M2_1440_420 0 0.008f
c1559 net8_M2_1520_420 0 0.008f
r780 net8_M2_1520_420 net8_M2_1600_420 4.8
c1560 net8_M2_1520_420 0 0.008f
c1561 net8_M2_1600_420 0 0.008f
r781 net8_M2_1600_420 net8_M2_1680_420 4.8
c1562 net8_M2_1600_420 0 0.008f
c1563 net8_M2_1680_420 0 0.008f
r782 net8_M2_1680_420 net8_M2_1760_420 4.8
c1564 net8_M2_1680_420 0 0.008f
c1565 net8_M2_1760_420 0 0.008f
r783 net8_M2_1760_420 net8_M2_1840_420 4.8
c1566 net8_M2_1760_420 0 0.008f
c1567 net8_M2_1840_420 0 0.008f
r784 net8_M2_1840_420 net8_M2_1920_420 4.8
c1568 net8_M2_1840_420 0 0.008f
c1569 net8_M2_1920_420 0 0.008f
r785 net8_M2_1920_420 net8_M2_2000_420 4.8
c1570 net8_M2_1920_420 0 0.008f
c1571 net8_M2_2000_420 0 0.008f
r786 net8_M2_2000_420 net8_M2_2080_420 4.8
c1572 net8_M2_2000_420 0 0.008f
c1573 net8_M2_2080_420 0 0.008f
r787 net8_M2_2080_420 net8_M2_2160_420 4.8
c1574 net8_M2_2080_420 0 0.008f
c1575 net8_M2_2160_420 0 0.008f
r788 net8_M2_2160_420 net8_M2_2240_420 4.8
c1576 net8_M2_2160_420 0 0.008f
c1577 net8_M2_2240_420 0 0.008f
r789 net8_M2_2240_420 net8_M2_2320_420 4.8
c1578 net8_M2_2240_420 0 0.008f
c1579 net8_M2_2320_420 0 0.008f
r790 net8_M2_2320_420 net8_M2_2400_420 4.8
c1580 net8_M2_2320_420 0 0.008f
c1581 net8_M2_2400_420 0 0.008f
r791 net8_M2_2400_420 net8_M2_2480_420 4.8
c1582 net8_M2_2400_420 0 0.008f
c1583 net8_M2_2480_420 0 0.008f
r792 net8_M2_2480_420 net8_M2_2560_420 4.8
c1584 net8_M2_2480_420 0 0.008f
c1585 net8_M2_2560_420 0 0.008f
r793 net8_M2_2560_420 net8_M2_2640_420 4.8
c1586 net8_M2_2560_420 0 0.008f
c1587 net8_M2_2640_420 0 0.008f
r794 net8_M2_2640_420 net8_M2_2720_420 4.8
c1588 net8_M2_2640_420 0 0.008f
c1589 net8_M2_2720_420 0 0.008f
r795 net8_M2_2720_420 net8_M2_2800_420 4.8
c1590 net8_M2_2720_420 0 0.008f
c1591 net8_M2_2800_420 0 0.008f
r796 net8_M2_2800_420 net8_M2_2880_420 4.8
c1592 net8_M2_2800_420 0 0.008f
c1593 net8_M2_2880_420 0 0.008f
r797 net8_M2_2880_420 net8_M2_2960_420 4.8
c1594 net8_M2_2880_420 0 0.008f
c1595 net8_M2_2960_420 0 0.008f
r798 net8_M2_2960_420 net8_M2_3040_420 4.8
c1596 net8_M2_2960_420 0 0.008f
c1597 net8_M2_3040_420 0 0.008f
r799 net8_M2_3040_420 net8_M2_3120_420 4.8
c1598 net8_M2_3040_420 0 0.008f
c1599 net8_M2_3120_420 0 0.008f
r800 net8_M2_3120_420 net8_M2_3200_420 4.8
c1600 net8_M2_3120_420 0 0.008f
c1601 net8_M2_3200_420 0 0.008f
r801 net8_M2_3200_420 net8_M2_3280_420 4.8
c1602 net8_M2_3200_420 0 0.008f
c1603 net8_M2_3280_420 0 0.008f
r802 net8_M2_3280_420 net8_M2_3360_420 4.8
c1604 net8_M2_3280_420 0 0.008f
c1605 net8_M2_3360_420 0 0.008f
r803 net8_M2_3360_420 net8_M2_3440_420 4.8
c1606 net8_M2_3360_420 0 0.008f
c1607 net8_M2_3440_420 0 0.008f
r804 net8_M2_3440_420 net8_M2_3520_420 4.8
c1608 net8_M2_3440_420 0 0.008f
c1609 net8_M2_3520_420 0 0.008f
r805 net8_M2_3520_420 net8_M2_3600_420 4.8
c1610 net8_M2_3520_420 0 0.008f
c1611 net8_M2_3600_420 0 0.008f
r806 net8_M2_3600_420 net8_M2_3680_420 4.8
c1612 net8_M2_3600_420 0 0.008f
c1613 net8_M2_3680_420 0 0.008f
r807 net8_M2_3680_420 net8_M2_3760_420 4.8
c1614 net8_M2_3680_420 0 0.008f
c1615 net8_M2_3760_420 0 0.008f
r808 net8_M2_3760_420 net8_M2_3840_420 4.8
c1616 net8_M2_3760_420 0 0.008f
c1617 net8_M2_3840_420 0 0.008f
r809 net8_M2_3840_420 net8_M2_3920_420 4.8
c1618 net8_M2_3840_420 0 0.008f
c1619 net8_M2_3920_420 0 0.008f
r810 net8_M2_3920_420 net8_M2_3956_420 2.1599999999999997
c1620 net8_M2_3920_420 0 0.0036f
c1621 net8_M2_3956_420 0 0.0036f
r811 id_M2_364_504 id_M2_444_504 4.8
c1622 id_M2_364_504 0 0.008f
c1623 id_M2_444_504 0 0.008f
r812 id_M2_444_504 id_M2_524_504 4.8
c1624 id_M2_444_504 0 0.008f
c1625 id_M2_524_504 0 0.008f
r813 id_M2_524_504 id_M2_604_504 4.8
c1626 id_M2_524_504 0 0.008f
c1627 id_M2_604_504 0 0.008f
r814 id_M2_604_504 id_M2_684_504 4.8
c1628 id_M2_604_504 0 0.008f
c1629 id_M2_684_504 0 0.008f
r815 id_M2_684_504 id_M2_764_504 4.8
c1630 id_M2_684_504 0 0.008f
c1631 id_M2_764_504 0 0.008f
r816 id_M2_764_504 id_M2_844_504 4.8
c1632 id_M2_764_504 0 0.008f
c1633 id_M2_844_504 0 0.008f
r817 id_M2_844_504 id_M2_924_504 4.8
c1634 id_M2_844_504 0 0.008f
c1635 id_M2_924_504 0 0.008f
r818 id_M2_924_504 id_M2_1004_504 4.8
c1636 id_M2_924_504 0 0.008f
c1637 id_M2_1004_504 0 0.008f
r819 id_M2_1004_504 id_M2_1084_504 4.8
c1638 id_M2_1004_504 0 0.008f
c1639 id_M2_1084_504 0 0.008f
r820 id_M2_1084_504 id_M2_1164_504 4.8
c1640 id_M2_1084_504 0 0.008f
c1641 id_M2_1164_504 0 0.008f
r821 id_M2_1164_504 id_M2_1244_504 4.8
c1642 id_M2_1164_504 0 0.008f
c1643 id_M2_1244_504 0 0.008f
r822 id_M2_1244_504 id_M2_1324_504 4.8
c1644 id_M2_1244_504 0 0.008f
c1645 id_M2_1324_504 0 0.008f
r823 id_M2_1324_504 id_M2_1404_504 4.8
c1646 id_M2_1324_504 0 0.008f
c1647 id_M2_1404_504 0 0.008f
r824 id_M2_1404_504 id_M2_1484_504 4.8
c1648 id_M2_1404_504 0 0.008f
c1649 id_M2_1484_504 0 0.008f
r825 id_M2_1484_504 id_M2_1564_504 4.8
c1650 id_M2_1484_504 0 0.008f
c1651 id_M2_1564_504 0 0.008f
r826 id_M2_1564_504 id_M2_1644_504 4.8
c1652 id_M2_1564_504 0 0.008f
c1653 id_M2_1644_504 0 0.008f
r827 id_M2_1644_504 id_M2_1724_504 4.8
c1654 id_M2_1644_504 0 0.008f
c1655 id_M2_1724_504 0 0.008f
r828 id_M2_1724_504 id_M2_1804_504 4.8
c1656 id_M2_1724_504 0 0.008f
c1657 id_M2_1804_504 0 0.008f
r829 id_M2_1804_504 id_M2_1884_504 4.8
c1658 id_M2_1804_504 0 0.008f
c1659 id_M2_1884_504 0 0.008f
r830 id_M2_1884_504 id_M2_1964_504 4.8
c1660 id_M2_1884_504 0 0.008f
c1661 id_M2_1964_504 0 0.008f
r831 id_M2_1964_504 id_M2_2044_504 4.8
c1662 id_M2_1964_504 0 0.008f
c1663 id_M2_2044_504 0 0.008f
r832 id_M2_2044_504 id_M2_2124_504 4.8
c1664 id_M2_2044_504 0 0.008f
c1665 id_M2_2124_504 0 0.008f
r833 id_M2_2124_504 id_M2_2204_504 4.8
c1666 id_M2_2124_504 0 0.008f
c1667 id_M2_2204_504 0 0.008f
r834 id_M2_2204_504 id_M2_2284_504 4.8
c1668 id_M2_2204_504 0 0.008f
c1669 id_M2_2284_504 0 0.008f
r835 id_M2_2284_504 id_M2_2364_504 4.8
c1670 id_M2_2284_504 0 0.008f
c1671 id_M2_2364_504 0 0.008f
r836 id_M2_2364_504 id_M2_2444_504 4.8
c1672 id_M2_2364_504 0 0.008f
c1673 id_M2_2444_504 0 0.008f
r837 id_M2_2444_504 id_M2_2524_504 4.8
c1674 id_M2_2444_504 0 0.008f
c1675 id_M2_2524_504 0 0.008f
r838 id_M2_2524_504 id_M2_2604_504 4.8
c1676 id_M2_2524_504 0 0.008f
c1677 id_M2_2604_504 0 0.008f
r839 id_M2_2604_504 id_M2_2684_504 4.8
c1678 id_M2_2604_504 0 0.008f
c1679 id_M2_2684_504 0 0.008f
r840 id_M2_2684_504 id_M2_2764_504 4.8
c1680 id_M2_2684_504 0 0.008f
c1681 id_M2_2764_504 0 0.008f
r841 id_M2_2764_504 id_M2_2844_504 4.8
c1682 id_M2_2764_504 0 0.008f
c1683 id_M2_2844_504 0 0.008f
r842 id_M2_2844_504 id_M2_2924_504 4.8
c1684 id_M2_2844_504 0 0.008f
c1685 id_M2_2924_504 0 0.008f
r843 id_M2_2924_504 id_M2_3004_504 4.8
c1686 id_M2_2924_504 0 0.008f
c1687 id_M2_3004_504 0 0.008f
r844 id_M2_3004_504 id_M2_3040_504 2.1599999999999997
c1688 id_M2_3004_504 0 0.0036f
c1689 id_M2_3040_504 0 0.0036f
r845 id_M2_400_504 id_M2_480_504 4.8
c1690 id_M2_400_504 0 0.008f
c1691 id_M2_480_504 0 0.008f
r846 id_M2_480_504 id_M2_560_504 4.8
c1692 id_M2_480_504 0 0.008f
c1693 id_M2_560_504 0 0.008f
r847 id_M2_560_504 id_M2_640_504 4.8
c1694 id_M2_560_504 0 0.008f
c1695 id_M2_640_504 0 0.008f
r848 id_M2_640_504 id_M2_720_504 4.8
c1696 id_M2_640_504 0 0.008f
c1697 id_M2_720_504 0 0.008f
r849 id_M2_720_504 id_M2_800_504 4.8
c1698 id_M2_720_504 0 0.008f
c1699 id_M2_800_504 0 0.008f
r850 id_M2_800_504 id_M2_880_504 4.8
c1700 id_M2_800_504 0 0.008f
c1701 id_M2_880_504 0 0.008f
r851 id_M2_880_504 id_M2_960_504 4.8
c1702 id_M2_880_504 0 0.008f
c1703 id_M2_960_504 0 0.008f
r852 id_M2_960_504 id_M2_1040_504 4.8
c1704 id_M2_960_504 0 0.008f
c1705 id_M2_1040_504 0 0.008f
r853 id_M2_1040_504 id_M2_1076_504 2.1599999999999997
c1706 id_M2_1040_504 0 0.0036f
c1707 id_M2_1076_504 0 0.0036f
r854 vinn_M2_2204_504 vinn_M2_2284_504 4.8
c1708 vinn_M2_2204_504 0 0.008f
c1709 vinn_M2_2284_504 0 0.008f
r855 vinn_M2_2284_504 vinn_M2_2364_504 4.8
c1710 vinn_M2_2284_504 0 0.008f
c1711 vinn_M2_2364_504 0 0.008f
r856 vinn_M2_2364_504 vinn_M2_2444_504 4.8
c1712 vinn_M2_2364_504 0 0.008f
c1713 vinn_M2_2444_504 0 0.008f
r857 vinn_M2_2444_504 vinn_M2_2524_504 4.8
c1714 vinn_M2_2444_504 0 0.008f
c1715 vinn_M2_2524_504 0 0.008f
r858 vinn_M2_2524_504 vinn_M2_2604_504 4.8
c1716 vinn_M2_2524_504 0 0.008f
c1717 vinn_M2_2604_504 0 0.008f
r859 vinn_M2_2604_504 vinn_M2_2684_504 4.8
c1718 vinn_M2_2604_504 0 0.008f
c1719 vinn_M2_2684_504 0 0.008f
r860 vinn_M2_2684_504 vinn_M2_2764_504 4.8
c1720 vinn_M2_2684_504 0 0.008f
c1721 vinn_M2_2764_504 0 0.008f
r861 vinn_M2_2764_504 vinn_M2_2844_504 4.8
c1722 vinn_M2_2764_504 0 0.008f
c1723 vinn_M2_2844_504 0 0.008f
r862 vinn_M2_2844_504 vinn_M2_2924_504 4.8
c1724 vinn_M2_2844_504 0 0.008f
c1725 vinn_M2_2924_504 0 0.008f
r863 vinn_M2_2924_504 vinn_M2_3004_504 4.8
c1726 vinn_M2_2924_504 0 0.008f
c1727 vinn_M2_3004_504 0 0.008f
r864 vinn_M2_3004_504 vinn_M2_3040_504 2.1599999999999997
c1728 vinn_M2_3004_504 0 0.0036f
c1729 vinn_M2_3040_504 0 0.0036f
r865 vinn_M2_400_504 vinn_M2_480_504 4.8
c1730 vinn_M2_400_504 0 0.008f
c1731 vinn_M2_480_504 0 0.008f
r866 vinn_M2_480_504 vinn_M2_560_504 4.8
c1732 vinn_M2_480_504 0 0.008f
c1733 vinn_M2_560_504 0 0.008f
r867 vinn_M2_560_504 vinn_M2_640_504 4.8
c1734 vinn_M2_560_504 0 0.008f
c1735 vinn_M2_640_504 0 0.008f
r868 vinn_M2_640_504 vinn_M2_720_504 4.8
c1736 vinn_M2_640_504 0 0.008f
c1737 vinn_M2_720_504 0 0.008f
r869 vinn_M2_720_504 vinn_M2_800_504 4.8
c1738 vinn_M2_720_504 0 0.008f
c1739 vinn_M2_800_504 0 0.008f
r870 vinn_M2_800_504 vinn_M2_880_504 4.8
c1740 vinn_M2_800_504 0 0.008f
c1741 vinn_M2_880_504 0 0.008f
r871 vinn_M2_880_504 vinn_M2_960_504 4.8
c1742 vinn_M2_880_504 0 0.008f
c1743 vinn_M2_960_504 0 0.008f
r872 vinn_M2_960_504 vinn_M2_1040_504 4.8
c1744 vinn_M2_960_504 0 0.008f
c1745 vinn_M2_1040_504 0 0.008f
r873 vinn_M2_1040_504 vinn_M2_1120_504 4.8
c1746 vinn_M2_1040_504 0 0.008f
c1747 vinn_M2_1120_504 0 0.008f
r874 vinn_M2_1120_504 vinn_M2_1200_504 4.8
c1748 vinn_M2_1120_504 0 0.008f
c1749 vinn_M2_1200_504 0 0.008f
r875 vinn_M2_1200_504 vinn_M2_1280_504 4.8
c1750 vinn_M2_1200_504 0 0.008f
c1751 vinn_M2_1280_504 0 0.008f
r876 vinn_M2_1280_504 vinn_M2_1360_504 4.8
c1752 vinn_M2_1280_504 0 0.008f
c1753 vinn_M2_1360_504 0 0.008f
r877 vinn_M2_1360_504 vinn_M2_1440_504 4.8
c1754 vinn_M2_1360_504 0 0.008f
c1755 vinn_M2_1440_504 0 0.008f
r878 vinn_M2_1440_504 vinn_M2_1520_504 4.8
c1756 vinn_M2_1440_504 0 0.008f
c1757 vinn_M2_1520_504 0 0.008f
r879 vinn_M2_1520_504 vinn_M2_1600_504 4.8
c1758 vinn_M2_1520_504 0 0.008f
c1759 vinn_M2_1600_504 0 0.008f
r880 vinn_M2_1600_504 vinn_M2_1680_504 4.8
c1760 vinn_M2_1600_504 0 0.008f
c1761 vinn_M2_1680_504 0 0.008f
r881 vinn_M2_1680_504 vinn_M2_1760_504 4.8
c1762 vinn_M2_1680_504 0 0.008f
c1763 vinn_M2_1760_504 0 0.008f
r882 vinn_M2_1760_504 vinn_M2_1840_504 4.8
c1764 vinn_M2_1760_504 0 0.008f
c1765 vinn_M2_1840_504 0 0.008f
r883 vinn_M2_1840_504 vinn_M2_1920_504 4.8
c1766 vinn_M2_1840_504 0 0.008f
c1767 vinn_M2_1920_504 0 0.008f
r884 vinn_M2_1920_504 vinn_M2_2000_504 4.8
c1768 vinn_M2_1920_504 0 0.008f
c1769 vinn_M2_2000_504 0 0.008f
r885 vinn_M2_2000_504 vinn_M2_2080_504 4.8
c1770 vinn_M2_2000_504 0 0.008f
c1771 vinn_M2_2080_504 0 0.008f
r886 vinn_M2_2080_504 vinn_M2_2160_504 4.8
c1772 vinn_M2_2080_504 0 0.008f
c1773 vinn_M2_2160_504 0 0.008f
r887 vinn_M2_2160_504 vinn_M2_2240_504 4.8
c1774 vinn_M2_2160_504 0 0.008f
c1775 vinn_M2_2240_504 0 0.008f
r888 vinn_M2_2240_504 vinn_M2_2320_504 4.8
c1776 vinn_M2_2240_504 0 0.008f
c1777 vinn_M2_2320_504 0 0.008f
r889 vinn_M2_2320_504 vinn_M2_2400_504 4.8
c1778 vinn_M2_2320_504 0 0.008f
c1779 vinn_M2_2400_504 0 0.008f
r890 vinn_M2_2400_504 vinn_M2_2436_504 2.1599999999999997
c1780 vinn_M2_2400_504 0 0.0036f
c1781 vinn_M2_2436_504 0 0.0036f
r891 vout_M2_2924_504 vout_M2_3004_504 4.8
c1782 vout_M2_2924_504 0 0.008f
c1783 vout_M2_3004_504 0 0.008f
r892 vout_M2_3004_504 vout_M2_3040_504 2.1599999999999997
c1784 vout_M2_3004_504 0 0.0036f
c1785 vout_M2_3040_504 0 0.0036f
r893 vout_M2_400_504 vout_M2_480_504 4.8
c1786 vout_M2_400_504 0 0.008f
c1787 vout_M2_480_504 0 0.008f
r894 vout_M2_480_504 vout_M2_560_504 4.8
c1788 vout_M2_480_504 0 0.008f
c1789 vout_M2_560_504 0 0.008f
r895 vout_M2_560_504 vout_M2_640_504 4.8
c1790 vout_M2_560_504 0 0.008f
c1791 vout_M2_640_504 0 0.008f
r896 vout_M2_640_504 vout_M2_720_504 4.8
c1792 vout_M2_640_504 0 0.008f
c1793 vout_M2_720_504 0 0.008f
r897 vout_M2_720_504 vout_M2_800_504 4.8
c1794 vout_M2_720_504 0 0.008f
c1795 vout_M2_800_504 0 0.008f
r898 vout_M2_800_504 vout_M2_880_504 4.8
c1796 vout_M2_800_504 0 0.008f
c1797 vout_M2_880_504 0 0.008f
r899 vout_M2_880_504 vout_M2_960_504 4.8
c1798 vout_M2_880_504 0 0.008f
c1799 vout_M2_960_504 0 0.008f
r900 vout_M2_960_504 vout_M2_1040_504 4.8
c1800 vout_M2_960_504 0 0.008f
c1801 vout_M2_1040_504 0 0.008f
r901 vout_M2_1040_504 vout_M2_1120_504 4.8
c1802 vout_M2_1040_504 0 0.008f
c1803 vout_M2_1120_504 0 0.008f
r902 vout_M2_1120_504 vout_M2_1200_504 4.8
c1804 vout_M2_1120_504 0 0.008f
c1805 vout_M2_1200_504 0 0.008f
r903 vout_M2_1200_504 vout_M2_1280_504 4.8
c1806 vout_M2_1200_504 0 0.008f
c1807 vout_M2_1280_504 0 0.008f
r904 vout_M2_1280_504 vout_M2_1360_504 4.8
c1808 vout_M2_1280_504 0 0.008f
c1809 vout_M2_1360_504 0 0.008f
r905 vout_M2_1360_504 vout_M2_1440_504 4.8
c1810 vout_M2_1360_504 0 0.008f
c1811 vout_M2_1440_504 0 0.008f
r906 vout_M2_1440_504 vout_M2_1520_504 4.8
c1812 vout_M2_1440_504 0 0.008f
c1813 vout_M2_1520_504 0 0.008f
r907 vout_M2_1520_504 vout_M2_1600_504 4.8
c1814 vout_M2_1520_504 0 0.008f
c1815 vout_M2_1600_504 0 0.008f
r908 vout_M2_1600_504 vout_M2_1680_504 4.8
c1816 vout_M2_1600_504 0 0.008f
c1817 vout_M2_1680_504 0 0.008f
r909 vout_M2_1680_504 vout_M2_1760_504 4.8
c1818 vout_M2_1680_504 0 0.008f
c1819 vout_M2_1760_504 0 0.008f
r910 vout_M2_1760_504 vout_M2_1840_504 4.8
c1820 vout_M2_1760_504 0 0.008f
c1821 vout_M2_1840_504 0 0.008f
r911 vout_M2_1840_504 vout_M2_1920_504 4.8
c1822 vout_M2_1840_504 0 0.008f
c1823 vout_M2_1920_504 0 0.008f
r912 vout_M2_1920_504 vout_M2_2000_504 4.8
c1824 vout_M2_1920_504 0 0.008f
c1825 vout_M2_2000_504 0 0.008f
r913 vout_M2_2000_504 vout_M2_2080_504 4.8
c1826 vout_M2_2000_504 0 0.008f
c1827 vout_M2_2080_504 0 0.008f
r914 vout_M2_2080_504 vout_M2_2160_504 4.8
c1828 vout_M2_2080_504 0 0.008f
c1829 vout_M2_2160_504 0 0.008f
r915 vout_M2_2160_504 vout_M2_2240_504 4.8
c1830 vout_M2_2160_504 0 0.008f
c1831 vout_M2_2240_504 0 0.008f
r916 vout_M2_2240_504 vout_M2_2320_504 4.8
c1832 vout_M2_2240_504 0 0.008f
c1833 vout_M2_2320_504 0 0.008f
r917 vout_M2_2320_504 vout_M2_2400_504 4.8
c1834 vout_M2_2320_504 0 0.008f
c1835 vout_M2_2400_504 0 0.008f
r918 vout_M2_2400_504 vout_M2_2480_504 4.8
c1836 vout_M2_2400_504 0 0.008f
c1837 vout_M2_2480_504 0 0.008f
r919 vout_M2_2480_504 vout_M2_2560_504 4.8
c1838 vout_M2_2480_504 0 0.008f
c1839 vout_M2_2560_504 0 0.008f
r920 vout_M2_2560_504 vout_M2_2640_504 4.8
c1840 vout_M2_2560_504 0 0.008f
c1841 vout_M2_2640_504 0 0.008f
r921 vout_M2_2640_504 vout_M2_2720_504 4.8
c1842 vout_M2_2640_504 0 0.008f
c1843 vout_M2_2720_504 0 0.008f
r922 vout_M2_2720_504 vout_M2_2800_504 4.8
c1844 vout_M2_2720_504 0 0.008f
c1845 vout_M2_2800_504 0 0.008f
r923 vout_M2_2800_504 vout_M2_2880_504 4.8
c1846 vout_M2_2800_504 0 0.008f
c1847 vout_M2_2880_504 0 0.008f
r924 vout_M2_2880_504 vout_M2_2960_504 4.8
c1848 vout_M2_2880_504 0 0.008f
c1849 vout_M2_2960_504 0 0.008f
r925 vout_M2_2960_504 vout_M2_3040_504 4.8
c1850 vout_M2_2960_504 0 0.008f
c1851 vout_M2_3040_504 0 0.008f
r926 vout_M2_3040_504 vout_M2_3120_504 4.8
c1852 vout_M2_3040_504 0 0.008f
c1853 vout_M2_3120_504 0 0.008f
r927 vout_M2_3120_504 vout_M2_3200_504 4.8
c1854 vout_M2_3120_504 0 0.008f
c1855 vout_M2_3200_504 0 0.008f
r928 vout_M2_3200_504 vout_M2_3236_504 2.1599999999999997
c1856 vout_M2_3200_504 0 0.0036f
c1857 vout_M2_3236_504 0 0.0036f
r929 net10_M2_684_588 net10_M2_764_588 4.8
c1858 net10_M2_684_588 0 0.008f
c1859 net10_M2_764_588 0 0.008f
r930 net10_M2_764_588 net10_M2_844_588 4.8
c1860 net10_M2_764_588 0 0.008f
c1861 net10_M2_844_588 0 0.008f
r931 net10_M2_844_588 net10_M2_924_588 4.8
c1862 net10_M2_844_588 0 0.008f
c1863 net10_M2_924_588 0 0.008f
r932 net10_M2_924_588 net10_M2_1004_588 4.8
c1864 net10_M2_924_588 0 0.008f
c1865 net10_M2_1004_588 0 0.008f
r933 net10_M2_1004_588 net10_M2_1084_588 4.8
c1866 net10_M2_1004_588 0 0.008f
c1867 net10_M2_1084_588 0 0.008f
r934 net10_M2_1084_588 net10_M2_1164_588 4.8
c1868 net10_M2_1084_588 0 0.008f
c1869 net10_M2_1164_588 0 0.008f
r935 net10_M2_1164_588 net10_M2_1244_588 4.8
c1870 net10_M2_1164_588 0 0.008f
c1871 net10_M2_1244_588 0 0.008f
r936 net10_M2_1244_588 net10_M2_1324_588 4.8
c1872 net10_M2_1244_588 0 0.008f
c1873 net10_M2_1324_588 0 0.008f
r937 net10_M2_1324_588 net10_M2_1404_588 4.8
c1874 net10_M2_1324_588 0 0.008f
c1875 net10_M2_1404_588 0 0.008f
r938 net10_M2_1404_588 net10_M2_1484_588 4.8
c1876 net10_M2_1404_588 0 0.008f
c1877 net10_M2_1484_588 0 0.008f
r939 net10_M2_1484_588 net10_M2_1564_588 4.8
c1878 net10_M2_1484_588 0 0.008f
c1879 net10_M2_1564_588 0 0.008f
r940 net10_M2_1564_588 net10_M2_1644_588 4.8
c1880 net10_M2_1564_588 0 0.008f
c1881 net10_M2_1644_588 0 0.008f
r941 net10_M2_1644_588 net10_M2_1724_588 4.8
c1882 net10_M2_1644_588 0 0.008f
c1883 net10_M2_1724_588 0 0.008f
r942 net10_M2_1724_588 net10_M2_1804_588 4.8
c1884 net10_M2_1724_588 0 0.008f
c1885 net10_M2_1804_588 0 0.008f
r943 net10_M2_1804_588 net10_M2_1884_588 4.8
c1886 net10_M2_1804_588 0 0.008f
c1887 net10_M2_1884_588 0 0.008f
r944 net10_M2_1884_588 net10_M2_1964_588 4.8
c1888 net10_M2_1884_588 0 0.008f
c1889 net10_M2_1964_588 0 0.008f
r945 net10_M2_1964_588 net10_M2_2044_588 4.8
c1890 net10_M2_1964_588 0 0.008f
c1891 net10_M2_2044_588 0 0.008f
r946 net10_M2_2044_588 net10_M2_2124_588 4.8
c1892 net10_M2_2044_588 0 0.008f
c1893 net10_M2_2124_588 0 0.008f
r947 net10_M2_2124_588 net10_M2_2204_588 4.8
c1894 net10_M2_2124_588 0 0.008f
c1895 net10_M2_2204_588 0 0.008f
r948 net10_M2_2204_588 net10_M2_2284_588 4.8
c1896 net10_M2_2204_588 0 0.008f
c1897 net10_M2_2284_588 0 0.008f
r949 net10_M2_2284_588 net10_M2_2364_588 4.8
c1898 net10_M2_2284_588 0 0.008f
c1899 net10_M2_2364_588 0 0.008f
r950 net10_M2_2364_588 net10_M2_2444_588 4.8
c1900 net10_M2_2364_588 0 0.008f
c1901 net10_M2_2444_588 0 0.008f
r951 net10_M2_2444_588 net10_M2_2524_588 4.8
c1902 net10_M2_2444_588 0 0.008f
c1903 net10_M2_2524_588 0 0.008f
r952 net10_M2_2524_588 net10_M2_2604_588 4.8
c1904 net10_M2_2524_588 0 0.008f
c1905 net10_M2_2604_588 0 0.008f
r953 net10_M2_2604_588 net10_M2_2684_588 4.8
c1906 net10_M2_2604_588 0 0.008f
c1907 net10_M2_2684_588 0 0.008f
r954 net10_M2_2684_588 net10_M2_2764_588 4.8
c1908 net10_M2_2684_588 0 0.008f
c1909 net10_M2_2764_588 0 0.008f
r955 net10_M2_2764_588 net10_M2_2844_588 4.8
c1910 net10_M2_2764_588 0 0.008f
c1911 net10_M2_2844_588 0 0.008f
r956 net10_M2_2844_588 net10_M2_2924_588 4.8
c1912 net10_M2_2844_588 0 0.008f
c1913 net10_M2_2924_588 0 0.008f
r957 net10_M2_2924_588 net10_M2_3004_588 4.8
c1914 net10_M2_2924_588 0 0.008f
c1915 net10_M2_3004_588 0 0.008f
r958 net10_M2_3004_588 net10_M2_3084_588 4.8
c1916 net10_M2_3004_588 0 0.008f
c1917 net10_M2_3084_588 0 0.008f
r959 net10_M2_3084_588 net10_M2_3120_588 2.1599999999999997
c1918 net10_M2_3084_588 0 0.0036f
c1919 net10_M2_3120_588 0 0.0036f
r960 net10_M2_1120_588 net10_M2_1156_588 2.1599999999999997
c1920 net10_M2_1120_588 0 0.0036f
c1921 net10_M2_1156_588 0 0.0036f
r961 net8_M2_2844_588 net8_M2_2924_588 4.8
c1922 net8_M2_2844_588 0 0.008f
c1923 net8_M2_2924_588 0 0.008f
r962 net8_M2_2924_588 net8_M2_3004_588 4.8
c1924 net8_M2_2924_588 0 0.008f
c1925 net8_M2_3004_588 0 0.008f
r963 net8_M2_3004_588 net8_M2_3084_588 4.8
c1926 net8_M2_3004_588 0 0.008f
c1927 net8_M2_3084_588 0 0.008f
r964 net8_M2_3084_588 net8_M2_3120_588 2.1599999999999997
c1928 net8_M2_3084_588 0 0.0036f
c1929 net8_M2_3120_588 0 0.0036f
r965 net8_M2_1120_588 net8_M2_1200_588 4.8
c1930 net8_M2_1120_588 0 0.008f
c1931 net8_M2_1200_588 0 0.008f
r966 net8_M2_1200_588 net8_M2_1280_588 4.8
c1932 net8_M2_1200_588 0 0.008f
c1933 net8_M2_1280_588 0 0.008f
r967 net8_M2_1280_588 net8_M2_1360_588 4.8
c1934 net8_M2_1280_588 0 0.008f
c1935 net8_M2_1360_588 0 0.008f
r968 net8_M2_1360_588 net8_M2_1440_588 4.8
c1936 net8_M2_1360_588 0 0.008f
c1937 net8_M2_1440_588 0 0.008f
r969 net8_M2_1440_588 net8_M2_1520_588 4.8
c1938 net8_M2_1440_588 0 0.008f
c1939 net8_M2_1520_588 0 0.008f
r970 net8_M2_1520_588 net8_M2_1600_588 4.8
c1940 net8_M2_1520_588 0 0.008f
c1941 net8_M2_1600_588 0 0.008f
r971 net8_M2_1600_588 net8_M2_1680_588 4.8
c1942 net8_M2_1600_588 0 0.008f
c1943 net8_M2_1680_588 0 0.008f
r972 net8_M2_1680_588 net8_M2_1760_588 4.8
c1944 net8_M2_1680_588 0 0.008f
c1945 net8_M2_1760_588 0 0.008f
r973 net8_M2_1760_588 net8_M2_1840_588 4.8
c1946 net8_M2_1760_588 0 0.008f
c1947 net8_M2_1840_588 0 0.008f
r974 net8_M2_1840_588 net8_M2_1920_588 4.8
c1948 net8_M2_1840_588 0 0.008f
c1949 net8_M2_1920_588 0 0.008f
r975 net8_M2_1920_588 net8_M2_2000_588 4.8
c1950 net8_M2_1920_588 0 0.008f
c1951 net8_M2_2000_588 0 0.008f
r976 net8_M2_2000_588 net8_M2_2080_588 4.8
c1952 net8_M2_2000_588 0 0.008f
c1953 net8_M2_2080_588 0 0.008f
r977 net8_M2_2080_588 net8_M2_2160_588 4.8
c1954 net8_M2_2080_588 0 0.008f
c1955 net8_M2_2160_588 0 0.008f
r978 net8_M2_2160_588 net8_M2_2240_588 4.8
c1956 net8_M2_2160_588 0 0.008f
c1957 net8_M2_2240_588 0 0.008f
r979 net8_M2_2240_588 net8_M2_2320_588 4.8
c1958 net8_M2_2240_588 0 0.008f
c1959 net8_M2_2320_588 0 0.008f
r980 net8_M2_2320_588 net8_M2_2400_588 4.8
c1960 net8_M2_2320_588 0 0.008f
c1961 net8_M2_2400_588 0 0.008f
r981 net8_M2_2400_588 net8_M2_2480_588 4.8
c1962 net8_M2_2400_588 0 0.008f
c1963 net8_M2_2480_588 0 0.008f
r982 net8_M2_2480_588 net8_M2_2560_588 4.8
c1964 net8_M2_2480_588 0 0.008f
c1965 net8_M2_2560_588 0 0.008f
r983 net8_M2_2560_588 net8_M2_2640_588 4.8
c1966 net8_M2_2560_588 0 0.008f
c1967 net8_M2_2640_588 0 0.008f
r984 net8_M2_2640_588 net8_M2_2720_588 4.8
c1968 net8_M2_2640_588 0 0.008f
c1969 net8_M2_2720_588 0 0.008f
r985 net8_M2_2720_588 net8_M2_2800_588 4.8
c1970 net8_M2_2720_588 0 0.008f
c1971 net8_M2_2800_588 0 0.008f
r986 net8_M2_2800_588 net8_M2_2880_588 4.8
c1972 net8_M2_2800_588 0 0.008f
c1973 net8_M2_2880_588 0 0.008f
r987 net8_M2_720_588 net8_M2_800_588 4.8
c1974 net8_M2_720_588 0 0.008f
c1975 net8_M2_800_588 0 0.008f
r988 net8_M2_800_588 net8_M2_880_588 4.8
c1976 net8_M2_800_588 0 0.008f
c1977 net8_M2_880_588 0 0.008f
r989 net8_M2_880_588 net8_M2_960_588 4.8
c1978 net8_M2_880_588 0 0.008f
c1979 net8_M2_960_588 0 0.008f
r990 net8_M2_960_588 net8_M2_1040_588 4.8
c1980 net8_M2_960_588 0 0.008f
c1981 net8_M2_1040_588 0 0.008f
r991 net8_M2_1040_588 net8_M2_1120_588 4.8
c1982 net8_M2_1040_588 0 0.008f
c1983 net8_M2_1120_588 0 0.008f
r992 net8_M2_2880_588 net8_M2_2960_588 4.8
c1984 net8_M2_2880_588 0 0.008f
c1985 net8_M2_2960_588 0 0.008f
r993 net8_M2_2960_588 net8_M2_3040_588 4.8
c1986 net8_M2_2960_588 0 0.008f
c1987 net8_M2_3040_588 0 0.008f
r994 net8_M2_3040_588 net8_M2_3120_588 4.8
c1988 net8_M2_3040_588 0 0.008f
c1989 net8_M2_3120_588 0 0.008f
r995 net8_M2_3120_588 net8_M2_3200_588 4.8
c1990 net8_M2_3120_588 0 0.008f
c1991 net8_M2_3200_588 0 0.008f
r996 net8_M2_3200_588 net8_M2_3236_588 2.1599999999999997
c1992 net8_M2_3200_588 0 0.0036f
c1993 net8_M2_3236_588 0 0.0036f
r997 id_M2_540_0 id_M2_620_0 4.8
c1994 id_M2_540_0 0 0.008f
c1995 id_M2_620_0 0 0.008f
r998 id_M2_620_0 id_M2_700_0 4.8
c1996 id_M2_620_0 0 0.008f
c1997 id_M2_700_0 0 0.008f
r999 id_M2_700_0 id_M2_780_0 4.8
c1998 id_M2_700_0 0 0.008f
c1999 id_M2_780_0 0 0.008f
r1000 id_M2_780_0 id_M2_860_0 4.8
c2000 id_M2_780_0 0 0.008f
c2001 id_M2_860_0 0 0.008f
r1001 id_M2_860_0 id_M2_940_0 4.8
c2002 id_M2_860_0 0 0.008f
c2003 id_M2_940_0 0 0.008f
r1002 id_M2_940_0 id_M2_1020_0 4.8
c2004 id_M2_940_0 0 0.008f
c2005 id_M2_1020_0 0 0.008f
r1003 id_M2_1020_0 id_M2_1100_0 4.8
c2006 id_M2_1020_0 0 0.008f
c2007 id_M2_1100_0 0 0.008f
r1004 id_M2_1100_0 id_M2_1180_0 4.8
c2008 id_M2_1100_0 0 0.008f
c2009 id_M2_1180_0 0 0.008f
r1005 id_M2_1180_0 id_M2_1260_0 4.8
c2010 id_M2_1180_0 0 0.008f
c2011 id_M2_1260_0 0 0.008f
r1006 id_M2_1260_0 id_M2_1340_0 4.8
c2012 id_M2_1260_0 0 0.008f
c2013 id_M2_1340_0 0 0.008f
r1007 id_M2_1340_0 id_M2_1420_0 4.8
c2014 id_M2_1340_0 0 0.008f
c2015 id_M2_1420_0 0 0.008f
r1008 id_M2_1420_0 id_M2_1500_0 4.8
c2016 id_M2_1420_0 0 0.008f
c2017 id_M2_1500_0 0 0.008f
r1009 id_M2_1500_0 id_M2_1580_0 4.8
c2018 id_M2_1500_0 0 0.008f
c2019 id_M2_1580_0 0 0.008f
r1010 id_M2_1580_0 id_M2_1660_0 4.8
c2020 id_M2_1580_0 0 0.008f
c2021 id_M2_1660_0 0 0.008f
r1011 id_M2_1660_0 id_M2_1740_0 4.8
c2022 id_M2_1660_0 0 0.008f
c2023 id_M2_1740_0 0 0.008f
r1012 id_M2_1740_0 id_M2_1820_0 4.8
c2024 id_M2_1740_0 0 0.008f
c2025 id_M2_1820_0 0 0.008f
r1013 id_M2_1820_0 id_M2_1900_0 4.8
c2026 id_M2_1820_0 0 0.008f
c2027 id_M2_1900_0 0 0.008f
r1014 id_M2_1900_0 id_M2_1980_0 4.8
c2028 id_M2_1900_0 0 0.008f
c2029 id_M2_1980_0 0 0.008f
r1015 id_M2_1980_0 id_M2_2060_0 4.8
c2030 id_M2_1980_0 0 0.008f
c2031 id_M2_2060_0 0 0.008f
r1016 id_M2_2060_0 id_M2_2140_0 4.8
c2032 id_M2_2060_0 0 0.008f
c2033 id_M2_2140_0 0 0.008f
r1017 id_M2_2140_0 id_M2_2220_0 4.8
c2034 id_M2_2140_0 0 0.008f
c2035 id_M2_2220_0 0 0.008f
r1018 id_M2_2220_0 id_M2_2300_0 4.8
c2036 id_M2_2220_0 0 0.008f
c2037 id_M2_2300_0 0 0.008f
r1019 id_M2_2300_0 id_M2_2380_0 4.8
c2038 id_M2_2300_0 0 0.008f
c2039 id_M2_2380_0 0 0.008f
r1020 id_M2_2380_0 id_M2_2460_0 4.8
c2040 id_M2_2380_0 0 0.008f
c2041 id_M2_2460_0 0 0.008f
r1021 id_M2_2460_0 id_M2_2540_0 4.8
c2042 id_M2_2460_0 0 0.008f
c2043 id_M2_2540_0 0 0.008f
r1022 id_M2_2540_0 id_M2_2620_0 4.8
c2044 id_M2_2540_0 0 0.008f
c2045 id_M2_2620_0 0 0.008f
r1023 id_M2_2620_0 id_M2_2700_0 4.8
c2046 id_M2_2620_0 0 0.008f
c2047 id_M2_2700_0 0 0.008f
r1024 id_M2_2700_0 id_M2_2780_0 4.8
c2048 id_M2_2700_0 0 0.008f
c2049 id_M2_2780_0 0 0.008f
r1025 id_M2_2780_0 id_M2_2860_0 4.8
c2050 id_M2_2780_0 0 0.008f
c2051 id_M2_2860_0 0 0.008f
r1026 id_M2_2860_0 id_M2_2940_0 4.8
c2052 id_M2_2860_0 0 0.008f
c2053 id_M2_2940_0 0 0.008f
r1027 id_M2_2940_0 id_M2_3020_0 4.8
c2054 id_M2_2940_0 0 0.008f
c2055 id_M2_3020_0 0 0.008f
r1028 id_M2_3020_0 id_M2_3100_0 4.8
c2056 id_M2_3020_0 0 0.008f
c2057 id_M2_3100_0 0 0.008f
r1029 id_M2_3100_0 id_M2_3180_0 4.8
c2058 id_M2_3100_0 0 0.008f
c2059 id_M2_3180_0 0 0.008f
r1030 id_M2_3180_0 id_M2_3260_0 4.8
c2060 id_M2_3180_0 0 0.008f
c2061 id_M2_3260_0 0 0.008f
r1031 id_M2_3260_0 id_M2_3340_0 4.8
c2062 id_M2_3260_0 0 0.008f
c2063 id_M2_3340_0 0 0.008f
r1032 id_M2_3340_0 id_M2_3420_0 4.8
c2064 id_M2_3340_0 0 0.008f
c2065 id_M2_3420_0 0 0.008f
r1033 id_M2_3420_0 id_M2_3500_0 4.8
c2066 id_M2_3420_0 0 0.008f
c2067 id_M2_3500_0 0 0.008f
r1034 id_M2_3500_0 id_M2_3580_0 4.8
c2068 id_M2_3500_0 0 0.008f
c2069 id_M2_3580_0 0 0.008f
r1035 id_M2_3580_0 id_M2_3660_0 4.8
c2070 id_M2_3580_0 0 0.008f
c2071 id_M2_3660_0 0 0.008f
r1036 id_M2_3660_0 id_M2_3740_0 4.8
c2072 id_M2_3660_0 0 0.008f
c2073 id_M2_3740_0 0 0.008f
r1037 id_M2_3740_0 id_M2_3820_0 4.8
c2074 id_M2_3740_0 0 0.008f
c2075 id_M2_3820_0 0 0.008f
r1038 id_M2_3820_0 id_M2_3900_0 4.8
c2076 id_M2_3820_0 0 0.008f
c2077 id_M2_3900_0 0 0.008f
r1039 id_M2_3900_0 id_M2_3920_0 1.2
c2078 id_M2_3900_0 0 0.002f
c2079 id_M2_3920_0 0 0.002f
r1040 id_M2_640_0 id_M2_720_0 4.8
c2080 id_M2_640_0 0 0.008f
c2081 id_M2_720_0 0 0.008f
r1041 id_M2_720_0 id_M2_740_0 1.2
c2082 id_M2_720_0 0 0.002f
c2083 id_M2_740_0 0 0.002f
r1042 vinp_M2_1324_0 vinp_M2_1404_0 4.8
c2084 vinp_M2_1324_0 0 0.008f
c2085 vinp_M2_1404_0 0 0.008f
r1043 vinp_M2_1404_0 vinp_M2_1484_0 4.8
c2086 vinp_M2_1404_0 0 0.008f
c2087 vinp_M2_1484_0 0 0.008f
r1044 vinp_M2_1484_0 vinp_M2_1564_0 4.8
c2088 vinp_M2_1484_0 0 0.008f
c2089 vinp_M2_1564_0 0 0.008f
r1045 vinp_M2_1564_0 vinp_M2_1644_0 4.8
c2090 vinp_M2_1564_0 0 0.008f
c2091 vinp_M2_1644_0 0 0.008f
r1046 vinp_M2_1644_0 vinp_M2_1724_0 4.8
c2092 vinp_M2_1644_0 0 0.008f
c2093 vinp_M2_1724_0 0 0.008f
r1047 vinp_M2_1724_0 vinp_M2_1804_0 4.8
c2094 vinp_M2_1724_0 0 0.008f
c2095 vinp_M2_1804_0 0 0.008f
r1048 vinp_M2_1804_0 vinp_M2_1884_0 4.8
c2096 vinp_M2_1804_0 0 0.008f
c2097 vinp_M2_1884_0 0 0.008f
r1049 vinp_M2_1884_0 vinp_M2_1964_0 4.8
c2098 vinp_M2_1884_0 0 0.008f
c2099 vinp_M2_1964_0 0 0.008f
r1050 vinp_M2_1964_0 vinp_M2_2044_0 4.8
c2100 vinp_M2_1964_0 0 0.008f
c2101 vinp_M2_2044_0 0 0.008f
r1051 vinp_M2_2044_0 vinp_M2_2124_0 4.8
c2102 vinp_M2_2044_0 0 0.008f
c2103 vinp_M2_2124_0 0 0.008f
r1052 vinp_M2_2124_0 vinp_M2_2204_0 4.8
c2104 vinp_M2_2124_0 0 0.008f
c2105 vinp_M2_2204_0 0 0.008f
r1053 vinp_M2_2204_0 vinp_M2_2284_0 4.8
c2106 vinp_M2_2204_0 0 0.008f
c2107 vinp_M2_2284_0 0 0.008f
r1054 vinp_M2_2284_0 vinp_M2_2364_0 4.8
c2108 vinp_M2_2284_0 0 0.008f
c2109 vinp_M2_2364_0 0 0.008f
r1055 vinp_M2_2364_0 vinp_M2_2444_0 4.8
c2110 vinp_M2_2364_0 0 0.008f
c2111 vinp_M2_2444_0 0 0.008f
r1056 vinp_M2_2444_0 vinp_M2_2524_0 4.8
c2112 vinp_M2_2444_0 0 0.008f
c2113 vinp_M2_2524_0 0 0.008f
r1057 vinp_M2_2524_0 vinp_M2_2604_0 4.8
c2114 vinp_M2_2524_0 0 0.008f
c2115 vinp_M2_2604_0 0 0.008f
r1058 vinp_M2_2604_0 vinp_M2_2684_0 4.8
c2116 vinp_M2_2604_0 0 0.008f
c2117 vinp_M2_2684_0 0 0.008f
r1059 vinp_M2_2684_0 vinp_M2_2764_0 4.8
c2118 vinp_M2_2684_0 0 0.008f
c2119 vinp_M2_2764_0 0 0.008f
r1060 vinp_M2_2764_0 vinp_M2_2844_0 4.8
c2120 vinp_M2_2764_0 0 0.008f
c2121 vinp_M2_2844_0 0 0.008f
r1061 vinp_M2_2844_0 vinp_M2_2924_0 4.8
c2122 vinp_M2_2844_0 0 0.008f
c2123 vinp_M2_2924_0 0 0.008f
r1062 vinp_M2_2924_0 vinp_M2_3004_0 4.8
c2124 vinp_M2_2924_0 0 0.008f
c2125 vinp_M2_3004_0 0 0.008f
r1063 vinp_M2_3004_0 vinp_M2_3084_0 4.8
c2126 vinp_M2_3004_0 0 0.008f
c2127 vinp_M2_3084_0 0 0.008f
r1064 vinp_M2_3084_0 vinp_M2_3164_0 4.8
c2128 vinp_M2_3084_0 0 0.008f
c2129 vinp_M2_3164_0 0 0.008f
r1065 vinp_M2_3164_0 vinp_M2_3244_0 4.8
c2130 vinp_M2_3164_0 0 0.008f
c2131 vinp_M2_3244_0 0 0.008f
r1066 vinp_M2_3244_0 vinp_M2_3324_0 4.8
c2132 vinp_M2_3244_0 0 0.008f
c2133 vinp_M2_3324_0 0 0.008f
r1067 vinp_M2_3324_0 vinp_M2_3404_0 4.8
c2134 vinp_M2_3324_0 0 0.008f
c2135 vinp_M2_3404_0 0 0.008f
r1068 vinp_M2_3404_0 vinp_M2_3484_0 4.8
c2136 vinp_M2_3404_0 0 0.008f
c2137 vinp_M2_3484_0 0 0.008f
r1069 vinp_M2_3484_0 vinp_M2_3564_0 4.8
c2138 vinp_M2_3484_0 0 0.008f
c2139 vinp_M2_3564_0 0 0.008f
r1070 vinp_M2_3564_0 vinp_M2_3644_0 4.8
c2140 vinp_M2_3564_0 0 0.008f
c2141 vinp_M2_3644_0 0 0.008f
r1071 vinp_M2_3644_0 vinp_M2_3724_0 4.8
c2142 vinp_M2_3644_0 0 0.008f
c2143 vinp_M2_3724_0 0 0.008f
r1072 vinp_M2_3724_0 vinp_M2_3804_0 4.8
c2144 vinp_M2_3724_0 0 0.008f
c2145 vinp_M2_3804_0 0 0.008f
r1073 vinp_M2_3804_0 vinp_M2_3884_0 4.8
c2146 vinp_M2_3804_0 0 0.008f
c2147 vinp_M2_3884_0 0 0.008f
r1074 vinp_M2_3884_0 vinp_M2_3920_0 2.1599999999999997
c2148 vinp_M2_3884_0 0 0.0036f
c2149 vinp_M2_3920_0 0 0.0036f
r1075 vinp_M2_640_0 vinp_M2_720_0 4.8
c2150 vinp_M2_640_0 0 0.008f
c2151 vinp_M2_720_0 0 0.008f
r1076 vinp_M2_720_0 vinp_M2_800_0 4.8
c2152 vinp_M2_720_0 0 0.008f
c2153 vinp_M2_800_0 0 0.008f
r1077 vinp_M2_800_0 vinp_M2_880_0 4.8
c2154 vinp_M2_800_0 0 0.008f
c2155 vinp_M2_880_0 0 0.008f
r1078 vinp_M2_880_0 vinp_M2_960_0 4.8
c2156 vinp_M2_880_0 0 0.008f
c2157 vinp_M2_960_0 0 0.008f
r1079 vinp_M2_960_0 vinp_M2_1040_0 4.8
c2158 vinp_M2_960_0 0 0.008f
c2159 vinp_M2_1040_0 0 0.008f
r1080 vinp_M2_1040_0 vinp_M2_1120_0 4.8
c2160 vinp_M2_1040_0 0 0.008f
c2161 vinp_M2_1120_0 0 0.008f
r1081 vinp_M2_1120_0 vinp_M2_1200_0 4.8
c2162 vinp_M2_1120_0 0 0.008f
c2163 vinp_M2_1200_0 0 0.008f
r1082 vinp_M2_1200_0 vinp_M2_1280_0 4.8
c2164 vinp_M2_1200_0 0 0.008f
c2165 vinp_M2_1280_0 0 0.008f
r1083 vinp_M2_1280_0 vinp_M2_1360_0 4.8
c2166 vinp_M2_1280_0 0 0.008f
c2167 vinp_M2_1360_0 0 0.008f
r1084 vinp_M2_1360_0 vinp_M2_1440_0 4.8
c2168 vinp_M2_1360_0 0 0.008f
c2169 vinp_M2_1440_0 0 0.008f
r1085 vinp_M2_1440_0 vinp_M2_1520_0 4.8
c2170 vinp_M2_1440_0 0 0.008f
c2171 vinp_M2_1520_0 0 0.008f
r1086 vinp_M2_1520_0 vinp_M2_1600_0 4.8
c2172 vinp_M2_1520_0 0 0.008f
c2173 vinp_M2_1600_0 0 0.008f
r1087 vinp_M2_1600_0 vinp_M2_1680_0 4.8
c2174 vinp_M2_1600_0 0 0.008f
c2175 vinp_M2_1680_0 0 0.008f
r1088 vinp_M2_1680_0 vinp_M2_1760_0 4.8
c2176 vinp_M2_1680_0 0 0.008f
c2177 vinp_M2_1760_0 0 0.008f
r1089 vinp_M2_1760_0 vinp_M2_1840_0 4.8
c2178 vinp_M2_1760_0 0 0.008f
c2179 vinp_M2_1840_0 0 0.008f
r1090 vout_M2_2300_0 vout_M2_2380_0 4.8
c2180 vout_M2_2300_0 0 0.008f
c2181 vout_M2_2380_0 0 0.008f
r1091 vout_M2_2380_0 vout_M2_2460_0 4.8
c2182 vout_M2_2380_0 0 0.008f
c2183 vout_M2_2460_0 0 0.008f
r1092 vout_M2_2460_0 vout_M2_2540_0 4.8
c2184 vout_M2_2460_0 0 0.008f
c2185 vout_M2_2540_0 0 0.008f
r1093 vout_M2_2540_0 vout_M2_2620_0 4.8
c2186 vout_M2_2540_0 0 0.008f
c2187 vout_M2_2620_0 0 0.008f
r1094 vout_M2_2620_0 vout_M2_2700_0 4.8
c2188 vout_M2_2620_0 0 0.008f
c2189 vout_M2_2700_0 0 0.008f
r1095 vout_M2_2700_0 vout_M2_2780_0 4.8
c2190 vout_M2_2700_0 0 0.008f
c2191 vout_M2_2780_0 0 0.008f
r1096 vout_M2_2780_0 vout_M2_2860_0 4.8
c2192 vout_M2_2780_0 0 0.008f
c2193 vout_M2_2860_0 0 0.008f
r1097 vout_M2_2860_0 vout_M2_2940_0 4.8
c2194 vout_M2_2860_0 0 0.008f
c2195 vout_M2_2940_0 0 0.008f
r1098 vout_M2_2940_0 vout_M2_3020_0 4.8
c2196 vout_M2_2940_0 0 0.008f
c2197 vout_M2_3020_0 0 0.008f
r1099 vout_M2_3020_0 vout_M2_3100_0 4.8
c2198 vout_M2_3020_0 0 0.008f
c2199 vout_M2_3100_0 0 0.008f
r1100 vout_M2_3100_0 vout_M2_3180_0 4.8
c2200 vout_M2_3100_0 0 0.008f
c2201 vout_M2_3180_0 0 0.008f
r1101 vout_M2_3180_0 vout_M2_3260_0 4.8
c2202 vout_M2_3180_0 0 0.008f
c2203 vout_M2_3260_0 0 0.008f
r1102 vout_M2_3260_0 vout_M2_3340_0 4.8
c2204 vout_M2_3260_0 0 0.008f
c2205 vout_M2_3340_0 0 0.008f
r1103 vout_M2_3340_0 vout_M2_3420_0 4.8
c2206 vout_M2_3340_0 0 0.008f
c2207 vout_M2_3420_0 0 0.008f
r1104 vout_M2_3420_0 vout_M2_3500_0 4.8
c2208 vout_M2_3420_0 0 0.008f
c2209 vout_M2_3500_0 0 0.008f
r1105 vout_M2_3500_0 vout_M2_3580_0 4.8
c2210 vout_M2_3500_0 0 0.008f
c2211 vout_M2_3580_0 0 0.008f
r1106 vout_M2_3580_0 vout_M2_3660_0 4.8
c2212 vout_M2_3580_0 0 0.008f
c2213 vout_M2_3660_0 0 0.008f
r1107 vout_M2_3660_0 vout_M2_3740_0 4.8
c2214 vout_M2_3660_0 0 0.008f
c2215 vout_M2_3740_0 0 0.008f
r1108 vout_M2_3740_0 vout_M2_3820_0 4.8
c2216 vout_M2_3740_0 0 0.008f
c2217 vout_M2_3820_0 0 0.008f
r1109 vout_M2_3820_0 vout_M2_3900_0 4.8
c2218 vout_M2_3820_0 0 0.008f
c2219 vout_M2_3900_0 0 0.008f
r1110 vout_M2_3900_0 vout_M2_3920_0 1.2
c2220 vout_M2_3900_0 0 0.002f
c2221 vout_M2_3920_0 0 0.002f
r1111 vout_M2_640_0 vout_M2_720_0 4.8
c2222 vout_M2_640_0 0 0.008f
c2223 vout_M2_720_0 0 0.008f
r1112 vout_M2_720_0 vout_M2_800_0 4.8
c2224 vout_M2_720_0 0 0.008f
c2225 vout_M2_800_0 0 0.008f
r1113 vout_M2_800_0 vout_M2_880_0 4.8
c2226 vout_M2_800_0 0 0.008f
c2227 vout_M2_880_0 0 0.008f
r1114 vout_M2_880_0 vout_M2_960_0 4.8
c2228 vout_M2_880_0 0 0.008f
c2229 vout_M2_960_0 0 0.008f
r1115 vout_M2_960_0 vout_M2_1040_0 4.8
c2230 vout_M2_960_0 0 0.008f
c2231 vout_M2_1040_0 0 0.008f
r1116 vout_M2_1040_0 vout_M2_1120_0 4.8
c2232 vout_M2_1040_0 0 0.008f
c2233 vout_M2_1120_0 0 0.008f
r1117 vout_M2_1120_0 vout_M2_1200_0 4.8
c2234 vout_M2_1120_0 0 0.008f
c2235 vout_M2_1200_0 0 0.008f
r1118 vout_M2_1200_0 vout_M2_1280_0 4.8
c2236 vout_M2_1200_0 0 0.008f
c2237 vout_M2_1280_0 0 0.008f
r1119 vout_M2_1280_0 vout_M2_1360_0 4.8
c2238 vout_M2_1280_0 0 0.008f
c2239 vout_M2_1360_0 0 0.008f
r1120 vout_M2_1360_0 vout_M2_1440_0 4.8
c2240 vout_M2_1360_0 0 0.008f
c2241 vout_M2_1440_0 0 0.008f
r1121 vout_M2_1440_0 vout_M2_1520_0 4.8
c2242 vout_M2_1440_0 0 0.008f
c2243 vout_M2_1520_0 0 0.008f
r1122 vout_M2_1520_0 vout_M2_1600_0 4.8
c2244 vout_M2_1520_0 0 0.008f
c2245 vout_M2_1600_0 0 0.008f
r1123 vout_M2_1600_0 vout_M2_1680_0 4.8
c2246 vout_M2_1600_0 0 0.008f
c2247 vout_M2_1680_0 0 0.008f
r1124 vout_M2_1680_0 vout_M2_1760_0 4.8
c2248 vout_M2_1680_0 0 0.008f
c2249 vout_M2_1760_0 0 0.008f
r1125 vout_M2_1760_0 vout_M2_1840_0 4.8
c2250 vout_M2_1760_0 0 0.008f
c2251 vout_M2_1840_0 0 0.008f
r1126 vout_M2_1840_0 vout_M2_1920_0 4.8
c2252 vout_M2_1840_0 0 0.008f
c2253 vout_M2_1920_0 0 0.008f
r1127 vout_M2_1920_0 vout_M2_2000_0 4.8
c2254 vout_M2_1920_0 0 0.008f
c2255 vout_M2_2000_0 0 0.008f
r1128 vout_M2_2000_0 vout_M2_2080_0 4.8
c2256 vout_M2_2000_0 0 0.008f
c2257 vout_M2_2080_0 0 0.008f
r1129 vout_M2_2080_0 vout_M2_2160_0 4.8
c2258 vout_M2_2080_0 0 0.008f
c2259 vout_M2_2160_0 0 0.008f
r1130 vout_M2_2160_0 vout_M2_2240_0 4.8
c2260 vout_M2_2160_0 0 0.008f
c2261 vout_M2_2240_0 0 0.008f
r1131 vout_M2_2240_0 vout_M2_2320_0 4.8
c2262 vout_M2_2240_0 0 0.008f
c2263 vout_M2_2320_0 0 0.008f
r1132 vout_M2_2320_0 vout_M2_2400_0 4.8
c2264 vout_M2_2320_0 0 0.008f
c2265 vout_M2_2400_0 0 0.008f
r1133 vout_M2_2400_0 vout_M2_2480_0 4.8
c2266 vout_M2_2400_0 0 0.008f
c2267 vout_M2_2480_0 0 0.008f
r1134 vout_M2_2480_0 vout_M2_2500_0 1.2
c2268 vout_M2_2480_0 0 0.002f
c2269 vout_M2_2500_0 0 0.002f
r1135 vdd_M2_3820_0 vdd_M2_3900_0 4.8
c2270 vdd_M2_3820_0 0 0.008f
c2271 vdd_M2_3900_0 0 0.008f
r1136 vdd_M2_3900_0 vdd_M2_3920_0 1.2
c2272 vdd_M2_3900_0 0 0.002f
c2273 vdd_M2_3920_0 0 0.002f
r1137 vdd_M2_640_0 vdd_M2_720_0 4.8
c2274 vdd_M2_640_0 0 0.008f
c2275 vdd_M2_720_0 0 0.008f
r1138 vdd_M2_720_0 vdd_M2_800_0 4.8
c2276 vdd_M2_720_0 0 0.008f
c2277 vdd_M2_800_0 0 0.008f
r1139 vdd_M2_800_0 vdd_M2_880_0 4.8
c2278 vdd_M2_800_0 0 0.008f
c2279 vdd_M2_880_0 0 0.008f
r1140 vdd_M2_880_0 vdd_M2_960_0 4.8
c2280 vdd_M2_880_0 0 0.008f
c2281 vdd_M2_960_0 0 0.008f
r1141 vdd_M2_960_0 vdd_M2_1040_0 4.8
c2282 vdd_M2_960_0 0 0.008f
c2283 vdd_M2_1040_0 0 0.008f
r1142 vdd_M2_1040_0 vdd_M2_1120_0 4.8
c2284 vdd_M2_1040_0 0 0.008f
c2285 vdd_M2_1120_0 0 0.008f
r1143 vdd_M2_1120_0 vdd_M2_1200_0 4.8
c2286 vdd_M2_1120_0 0 0.008f
c2287 vdd_M2_1200_0 0 0.008f
r1144 vdd_M2_1200_0 vdd_M2_1280_0 4.8
c2288 vdd_M2_1200_0 0 0.008f
c2289 vdd_M2_1280_0 0 0.008f
r1145 vdd_M2_1280_0 vdd_M2_1360_0 4.8
c2290 vdd_M2_1280_0 0 0.008f
c2291 vdd_M2_1360_0 0 0.008f
r1146 vdd_M2_1360_0 vdd_M2_1440_0 4.8
c2292 vdd_M2_1360_0 0 0.008f
c2293 vdd_M2_1440_0 0 0.008f
r1147 vdd_M2_1440_0 vdd_M2_1520_0 4.8
c2294 vdd_M2_1440_0 0 0.008f
c2295 vdd_M2_1520_0 0 0.008f
r1148 vdd_M2_1520_0 vdd_M2_1600_0 4.8
c2296 vdd_M2_1520_0 0 0.008f
c2297 vdd_M2_1600_0 0 0.008f
r1149 vdd_M2_1600_0 vdd_M2_1680_0 4.8
c2298 vdd_M2_1600_0 0 0.008f
c2299 vdd_M2_1680_0 0 0.008f
r1150 vdd_M2_1680_0 vdd_M2_1760_0 4.8
c2300 vdd_M2_1680_0 0 0.008f
c2301 vdd_M2_1760_0 0 0.008f
r1151 vdd_M2_1760_0 vdd_M2_1840_0 4.8
c2302 vdd_M2_1760_0 0 0.008f
c2303 vdd_M2_1840_0 0 0.008f
r1152 vdd_M2_1840_0 vdd_M2_1920_0 4.8
c2304 vdd_M2_1840_0 0 0.008f
c2305 vdd_M2_1920_0 0 0.008f
r1153 vdd_M2_1920_0 vdd_M2_2000_0 4.8
c2306 vdd_M2_1920_0 0 0.008f
c2307 vdd_M2_2000_0 0 0.008f
r1154 vdd_M2_2000_0 vdd_M2_2080_0 4.8
c2308 vdd_M2_2000_0 0 0.008f
c2309 vdd_M2_2080_0 0 0.008f
r1155 vdd_M2_2080_0 vdd_M2_2160_0 4.8
c2310 vdd_M2_2080_0 0 0.008f
c2311 vdd_M2_2160_0 0 0.008f
r1156 vdd_M2_2160_0 vdd_M2_2240_0 4.8
c2312 vdd_M2_2160_0 0 0.008f
c2313 vdd_M2_2240_0 0 0.008f
r1157 vdd_M2_2240_0 vdd_M2_2320_0 4.8
c2314 vdd_M2_2240_0 0 0.008f
c2315 vdd_M2_2320_0 0 0.008f
r1158 vdd_M2_2320_0 vdd_M2_2400_0 4.8
c2316 vdd_M2_2320_0 0 0.008f
c2317 vdd_M2_2400_0 0 0.008f
r1159 vdd_M2_2400_0 vdd_M2_2480_0 4.8
c2318 vdd_M2_2400_0 0 0.008f
c2319 vdd_M2_2480_0 0 0.008f
r1160 vdd_M2_2480_0 vdd_M2_2560_0 4.8
c2320 vdd_M2_2480_0 0 0.008f
c2321 vdd_M2_2560_0 0 0.008f
r1161 vdd_M2_2560_0 vdd_M2_2640_0 4.8
c2322 vdd_M2_2560_0 0 0.008f
c2323 vdd_M2_2640_0 0 0.008f
r1162 vdd_M2_2640_0 vdd_M2_2720_0 4.8
c2324 vdd_M2_2640_0 0 0.008f
c2325 vdd_M2_2720_0 0 0.008f
r1163 vdd_M2_2720_0 vdd_M2_2800_0 4.8
c2326 vdd_M2_2720_0 0 0.008f
c2327 vdd_M2_2800_0 0 0.008f
r1164 vdd_M2_2800_0 vdd_M2_2880_0 4.8
c2328 vdd_M2_2800_0 0 0.008f
c2329 vdd_M2_2880_0 0 0.008f
r1165 vdd_M2_2880_0 vdd_M2_2960_0 4.8
c2330 vdd_M2_2880_0 0 0.008f
c2331 vdd_M2_2960_0 0 0.008f
r1166 vdd_M2_2960_0 vdd_M2_3040_0 4.8
c2332 vdd_M2_2960_0 0 0.008f
c2333 vdd_M2_3040_0 0 0.008f
r1167 vdd_M2_3040_0 vdd_M2_3120_0 4.8
c2334 vdd_M2_3040_0 0 0.008f
c2335 vdd_M2_3120_0 0 0.008f
r1168 vdd_M2_3120_0 vdd_M2_3200_0 4.8
c2336 vdd_M2_3120_0 0 0.008f
c2337 vdd_M2_3200_0 0 0.008f
r1169 vdd_M2_3200_0 vdd_M2_3280_0 4.8
c2338 vdd_M2_3200_0 0 0.008f
c2339 vdd_M2_3280_0 0 0.008f
r1170 vdd_M2_3280_0 vdd_M2_3360_0 4.8
c2340 vdd_M2_3280_0 0 0.008f
c2341 vdd_M2_3360_0 0 0.008f
r1171 vdd_M2_3360_0 vdd_M2_3440_0 4.8
c2342 vdd_M2_3360_0 0 0.008f
c2343 vdd_M2_3440_0 0 0.008f
r1172 vdd_M2_3440_0 vdd_M2_3520_0 4.8
c2344 vdd_M2_3440_0 0 0.008f
c2345 vdd_M2_3520_0 0 0.008f
r1173 vdd_M2_3520_0 vdd_M2_3600_0 4.8
c2346 vdd_M2_3520_0 0 0.008f
c2347 vdd_M2_3600_0 0 0.008f
r1174 vdd_M2_3600_0 vdd_M2_3680_0 4.8
c2348 vdd_M2_3600_0 0 0.008f
c2349 vdd_M2_3680_0 0 0.008f
r1175 vdd_M2_3680_0 vdd_M2_3760_0 4.8
c2350 vdd_M2_3680_0 0 0.008f
c2351 vdd_M2_3760_0 0 0.008f
r1176 vdd_M2_3760_0 vdd_M2_3840_0 4.8
c2352 vdd_M2_3760_0 0 0.008f
c2353 vdd_M2_3840_0 0 0.008f
r1177 vdd_M2_3840_0 vdd_M2_3920_0 4.8
c2354 vdd_M2_3840_0 0 0.008f
c2355 vdd_M2_3920_0 0 0.008f
r1178 vdd_M2_3920_0 vdd_M2_4000_0 4.8
c2356 vdd_M2_3920_0 0 0.008f
c2357 vdd_M2_4000_0 0 0.008f
r1179 vdd_M2_4000_0 vdd_M2_4020_0 1.2
c2358 vdd_M2_4000_0 0 0.002f
c2359 vdd_M2_4020_0 0 0.002f
r1180 vout_M2_2444_84 vout_M2_2524_84 4.8
c2360 vout_M2_2444_84 0 0.008f
c2361 vout_M2_2524_84 0 0.008f
r1181 vout_M2_2524_84 vout_M2_2604_84 4.8
c2362 vout_M2_2524_84 0 0.008f
c2363 vout_M2_2604_84 0 0.008f
r1182 vout_M2_2604_84 vout_M2_2684_84 4.8
c2364 vout_M2_2604_84 0 0.008f
c2365 vout_M2_2684_84 0 0.008f
r1183 vout_M2_2684_84 vout_M2_2764_84 4.8
c2366 vout_M2_2684_84 0 0.008f
c2367 vout_M2_2764_84 0 0.008f
r1184 vout_M2_2764_84 vout_M2_2844_84 4.8
c2368 vout_M2_2764_84 0 0.008f
c2369 vout_M2_2844_84 0 0.008f
r1185 vout_M2_2844_84 vout_M2_2924_84 4.8
c2370 vout_M2_2844_84 0 0.008f
c2371 vout_M2_2924_84 0 0.008f
r1186 vout_M2_2924_84 vout_M2_2960_84 2.1599999999999997
c2372 vout_M2_2924_84 0 0.0036f
c2373 vout_M2_2960_84 0 0.0036f
r1187 vout_M2_2480_84 vout_M2_2560_84 4.8
c2374 vout_M2_2480_84 0 0.008f
c2375 vout_M2_2560_84 0 0.008f
r1188 vout_M2_2560_84 vout_M2_2640_84 4.8
c2376 vout_M2_2560_84 0 0.008f
c2377 vout_M2_2640_84 0 0.008f
r1189 vout_M2_2640_84 vout_M2_2720_84 4.8
c2378 vout_M2_2640_84 0 0.008f
c2379 vout_M2_2720_84 0 0.008f
r1190 vout_M2_2720_84 vout_M2_2800_84 4.8
c2380 vout_M2_2720_84 0 0.008f
c2381 vout_M2_2800_84 0 0.008f
r1191 vout_M2_2800_84 vout_M2_2880_84 4.8
c2382 vout_M2_2800_84 0 0.008f
c2383 vout_M2_2880_84 0 0.008f
r1192 vout_M2_2880_84 vout_M2_2960_84 4.8
c2384 vout_M2_2880_84 0 0.008f
c2385 vout_M2_2960_84 0 0.008f
r1193 vout_M2_2960_84 vout_M2_2996_84 2.1599999999999997
c2386 vout_M2_2960_84 0 0.0036f
c2387 vout_M2_2996_84 0 0.0036f
r1194 vdd_M1_3920_168 vdd_M2_3920_168 50
r1195 vdd_M1_3920_336 vdd_M2_3920_336 50
r1196 net8_M1_3840_252 net8_M2_3840_252 50
r1197 net8_M1_3840_420 net8_M2_3840_420 50
r1198 net8_M1_3760_252 net8_M2_3760_252 50
r1199 net8_M1_3760_420 net8_M2_3760_420 50
r1200 vdd_M1_3200_168 vdd_M2_3200_168 50
r1201 vdd_M1_3200_420 vdd_M2_3200_420 50
r1202 vout_M1_3040_252 vout_M2_3040_252 50
r1203 vout_M1_3040_504 vout_M2_3040_504 50
r1204 net8_M1_3120_336 net8_M2_3120_336 50
r1205 net8_M1_3120_588 net8_M2_3120_588 50
r1206 vss_M1_960_168 vss_M2_960_168 50
r1207 vss_M1_960_420 vss_M2_960_420 50
r1208 vss_M1_320_168 vss_M2_320_168 50
r1209 vss_M1_320_420 vss_M2_320_420 50
r1210 id_M1_1040_252 id_M2_1040_252 50
r1211 id_M1_1040_504 id_M2_1040_504 50
r1212 id_M1_400_252 id_M2_400_252 50
r1213 id_M1_400_504 id_M2_400_504 50
r1214 id_M1_480_252 id_M2_480_252 50
r1215 id_M1_480_504 id_M2_480_504 50
r1216 net10_M1_1120_336 net10_M2_1120_336 50
r1217 net10_M1_1120_588 net10_M2_1120_588 50
r1218 net10_M1_2320_168 net10_M2_2320_168 50
r1219 net10_M1_1680_168 net10_M2_1680_168 50
r1220 net8_M1_1840_252 net8_M2_1840_252 50
r1221 vout_M1_2480_336 vout_M2_2480_336 50
r1222 vinp_M1_1760_420 vinp_M2_1760_420 50
r1223 vinn_M1_2400_504 vinn_M2_2400_504 50
r1224 vdd_M3_3920__36 vdd_M3_3920_0 1.44
c2388 vdd_M3_3920__36 0 0.0036f
c2389 vdd_M3_3920_0 0 0.0036f
r1225 vdd_M3_3920_0 vdd_M3_3920_80 3.2
c2390 vdd_M3_3920_0 0 0.008f
c2391 vdd_M3_3920_80 0 0.008f
r1226 vdd_M3_3920_80 vdd_M3_3920_160 3.2
c2392 vdd_M3_3920_80 0 0.008f
c2393 vdd_M3_3920_160 0 0.008f
r1227 vdd_M3_3920_160 vdd_M3_3920_168 0.32
c2394 vdd_M3_3920_160 0 0.0008f
c2395 vdd_M3_3920_168 0 0.0008f
r1228 vdd_M3_3920_168 vdd_M3_3920_248 3.2
c2396 vdd_M3_3920_168 0 0.008f
c2397 vdd_M3_3920_248 0 0.008f
r1229 vdd_M3_3920_248 vdd_M3_3920_328 3.2
c2398 vdd_M3_3920_248 0 0.008f
c2399 vdd_M3_3920_328 0 0.008f
r1230 vdd_M3_3920_328 vdd_M3_3920_336 0.32
c2400 vdd_M3_3920_328 0 0.0008f
c2401 vdd_M3_3920_336 0 0.0008f
r1231 vdd_M3_3920_336 vdd_M3_3920_372 1.44
c2402 vdd_M3_3920_336 0 0.0036f
c2403 vdd_M3_3920_372 0 0.0036f
r1232 vdd_M3_3760_132 vdd_M3_3760_168 1.44
c2404 vdd_M3_3760_132 0 0.0036f
c2405 vdd_M3_3760_168 0 0.0036f
r1233 vdd_M3_3760_168 vdd_M3_3760_248 3.2
c2406 vdd_M3_3760_168 0 0.008f
c2407 vdd_M3_3760_248 0 0.008f
r1234 vdd_M3_3760_248 vdd_M3_3760_328 3.2
c2408 vdd_M3_3760_248 0 0.008f
c2409 vdd_M3_3760_328 0 0.008f
r1235 vdd_M3_3760_328 vdd_M3_3760_336 0.32
c2410 vdd_M3_3760_328 0 0.0008f
c2411 vdd_M3_3760_336 0 0.0008f
r1236 vdd_M3_3760_336 vdd_M3_3760_416 3.2
c2412 vdd_M3_3760_336 0 0.008f
c2413 vdd_M3_3760_416 0 0.008f
r1237 vdd_M3_3760_416 vdd_M3_3760_441 1.0
c2414 vdd_M3_3760_416 0 0.0025000000000000005f
c2415 vdd_M3_3760_441 0 0.0025000000000000005f
r1238 net8_M3_3840_216 net8_M3_3840_252 1.44
c2416 net8_M3_3840_216 0 0.0036f
c2417 net8_M3_3840_252 0 0.0036f
r1239 net8_M3_3840_252 net8_M3_3840_332 3.2
c2418 net8_M3_3840_252 0 0.008f
c2419 net8_M3_3840_332 0 0.008f
r1240 net8_M3_3840_332 net8_M3_3840_412 3.2
c2420 net8_M3_3840_332 0 0.008f
c2421 net8_M3_3840_412 0 0.008f
r1241 net8_M3_3840_412 net8_M3_3840_420 0.32
c2422 net8_M3_3840_412 0 0.0008f
c2423 net8_M3_3840_420 0 0.0008f
r1242 net8_M3_3840_420 net8_M3_3840_456 1.44
c2424 net8_M3_3840_420 0 0.0036f
c2425 net8_M3_3840_456 0 0.0036f
r1243 net8_M3_3680_216 net8_M3_3680_252 1.44
c2426 net8_M3_3680_216 0 0.0036f
c2427 net8_M3_3680_252 0 0.0036f
r1244 net8_M3_3680_252 net8_M3_3680_332 3.2
c2428 net8_M3_3680_252 0 0.008f
c2429 net8_M3_3680_332 0 0.008f
r1245 net8_M3_3680_332 net8_M3_3680_412 3.2
c2430 net8_M3_3680_332 0 0.008f
c2431 net8_M3_3680_412 0 0.008f
r1246 net8_M3_3680_412 net8_M3_3680_420 0.32
c2432 net8_M3_3680_412 0 0.0008f
c2433 net8_M3_3680_420 0 0.0008f
r1247 net8_M3_3680_420 net8_M3_3680_500 3.2
c2434 net8_M3_3680_420 0 0.008f
c2435 net8_M3_3680_500 0 0.008f
r1248 net8_M3_3680_500 net8_M3_3680_525 1.0
c2436 net8_M3_3680_500 0 0.0025000000000000005f
c2437 net8_M3_3680_525 0 0.0025000000000000005f
r1249 vdd_M3_3280_132 vdd_M3_3280_168 1.44
c2438 vdd_M3_3280_132 0 0.0036f
c2439 vdd_M3_3280_168 0 0.0036f
r1250 vdd_M3_3280_168 vdd_M3_3280_248 3.2
c2440 vdd_M3_3280_168 0 0.008f
c2441 vdd_M3_3280_248 0 0.008f
r1251 vdd_M3_3280_248 vdd_M3_3280_328 3.2
c2442 vdd_M3_3280_248 0 0.008f
c2443 vdd_M3_3280_328 0 0.008f
r1252 vdd_M3_3280_328 vdd_M3_3280_408 3.2
c2444 vdd_M3_3280_328 0 0.008f
c2445 vdd_M3_3280_408 0 0.008f
r1253 vdd_M3_3280_408 vdd_M3_3280_420 0.48
c2446 vdd_M3_3280_408 0 0.0012000000000000001f
c2447 vdd_M3_3280_420 0 0.0012000000000000001f
r1254 vdd_M3_3280_420 vdd_M3_3280_456 1.44
c2448 vdd_M3_3280_420 0 0.0036f
c2449 vdd_M3_3280_456 0 0.0036f
r1255 vdd_M3_3040_132 vdd_M3_3040_168 1.44
c2450 vdd_M3_3040_132 0 0.0036f
c2451 vdd_M3_3040_168 0 0.0036f
r1256 vdd_M3_3040_168 vdd_M3_3040_248 3.2
c2452 vdd_M3_3040_168 0 0.008f
c2453 vdd_M3_3040_248 0 0.008f
r1257 vdd_M3_3040_248 vdd_M3_3040_328 3.2
c2454 vdd_M3_3040_248 0 0.008f
c2455 vdd_M3_3040_328 0 0.008f
r1258 vdd_M3_3040_328 vdd_M3_3040_408 3.2
c2456 vdd_M3_3040_328 0 0.008f
c2457 vdd_M3_3040_408 0 0.008f
r1259 vdd_M3_3040_408 vdd_M3_3040_420 0.48
c2458 vdd_M3_3040_408 0 0.0012000000000000001f
c2459 vdd_M3_3040_420 0 0.0012000000000000001f
r1260 vdd_M3_3040_336 vdd_M3_3040_416 3.2
c2460 vdd_M3_3040_336 0 0.008f
c2461 vdd_M3_3040_416 0 0.008f
r1261 vdd_M3_3040_416 vdd_M3_3040_456 1.6
c2462 vdd_M3_3040_416 0 0.004f
c2463 vdd_M3_3040_456 0 0.004f
r1262 vout_M3_3200_216 vout_M3_3200_252 1.44
c2464 vout_M3_3200_216 0 0.0036f
c2465 vout_M3_3200_252 0 0.0036f
r1263 vout_M3_3200_252 vout_M3_3200_332 3.2
c2466 vout_M3_3200_252 0 0.008f
c2467 vout_M3_3200_332 0 0.008f
r1264 vout_M3_3200_332 vout_M3_3200_412 3.2
c2468 vout_M3_3200_332 0 0.008f
c2469 vout_M3_3200_412 0 0.008f
r1265 vout_M3_3200_412 vout_M3_3200_492 3.2
c2470 vout_M3_3200_412 0 0.008f
c2471 vout_M3_3200_492 0 0.008f
r1266 vout_M3_3200_492 vout_M3_3200_504 0.48
c2472 vout_M3_3200_492 0 0.0012000000000000001f
c2473 vout_M3_3200_504 0 0.0012000000000000001f
r1267 vout_M3_3200_504 vout_M3_3200_540 1.44
c2474 vout_M3_3200_504 0 0.0036f
c2475 vout_M3_3200_540 0 0.0036f
r1268 vout_M3_2960_48 vout_M3_2960_84 1.44
c2476 vout_M3_2960_48 0 0.0036f
c2477 vout_M3_2960_84 0 0.0036f
r1269 vout_M3_2960_84 vout_M3_2960_164 3.2
c2478 vout_M3_2960_84 0 0.008f
c2479 vout_M3_2960_164 0 0.008f
r1270 vout_M3_2960_164 vout_M3_2960_244 3.2
c2480 vout_M3_2960_164 0 0.008f
c2481 vout_M3_2960_244 0 0.008f
r1271 vout_M3_2960_244 vout_M3_2960_252 0.32
c2482 vout_M3_2960_244 0 0.0008f
c2483 vout_M3_2960_252 0 0.0008f
r1272 vout_M3_2960_252 vout_M3_2960_332 3.2
c2484 vout_M3_2960_252 0 0.008f
c2485 vout_M3_2960_332 0 0.008f
r1273 vout_M3_2960_332 vout_M3_2960_412 3.2
c2486 vout_M3_2960_332 0 0.008f
c2487 vout_M3_2960_412 0 0.008f
r1274 vout_M3_2960_412 vout_M3_2960_492 3.2
c2488 vout_M3_2960_412 0 0.008f
c2489 vout_M3_2960_492 0 0.008f
r1275 vout_M3_2960_492 vout_M3_2960_504 0.48
c2490 vout_M3_2960_492 0 0.0012000000000000001f
c2491 vout_M3_2960_504 0 0.0012000000000000001f
r1276 vout_M3_2960_504 vout_M3_2960_540 1.44
c2492 vout_M3_2960_504 0 0.0036f
c2493 vout_M3_2960_540 0 0.0036f
r1277 net8_M3_3120_300 net8_M3_3120_336 1.44
c2494 net8_M3_3120_300 0 0.0036f
c2495 net8_M3_3120_336 0 0.0036f
r1278 net8_M3_3120_336 net8_M3_3120_416 3.2
c2496 net8_M3_3120_336 0 0.008f
c2497 net8_M3_3120_416 0 0.008f
r1279 net8_M3_3120_416 net8_M3_3120_496 3.2
c2498 net8_M3_3120_416 0 0.008f
c2499 net8_M3_3120_496 0 0.008f
r1280 net8_M3_3120_496 net8_M3_3120_576 3.2
c2500 net8_M3_3120_496 0 0.008f
c2501 net8_M3_3120_576 0 0.008f
r1281 net8_M3_3120_576 net8_M3_3120_588 0.48
c2502 net8_M3_3120_576 0 0.0012000000000000001f
c2503 net8_M3_3120_588 0 0.0012000000000000001f
r1282 net8_M3_3120_588 net8_M3_3120_624 1.44
c2504 net8_M3_3120_588 0 0.0036f
c2505 net8_M3_3120_624 0 0.0036f
r1283 net8_M3_2880_300 net8_M3_2880_336 1.44
c2506 net8_M3_2880_300 0 0.0036f
c2507 net8_M3_2880_336 0 0.0036f
r1284 net8_M3_2880_336 net8_M3_2880_416 3.2
c2508 net8_M3_2880_336 0 0.008f
c2509 net8_M3_2880_416 0 0.008f
r1285 net8_M3_2880_416 net8_M3_2880_496 3.2
c2510 net8_M3_2880_416 0 0.008f
c2511 net8_M3_2880_496 0 0.008f
r1286 net8_M3_2880_496 net8_M3_2880_576 3.2
c2512 net8_M3_2880_496 0 0.008f
c2513 net8_M3_2880_576 0 0.008f
r1287 net8_M3_2880_576 net8_M3_2880_588 0.48
c2514 net8_M3_2880_576 0 0.0012000000000000001f
c2515 net8_M3_2880_588 0 0.0012000000000000001f
r1288 net8_M3_2880_420 net8_M3_2880_500 3.2
c2516 net8_M3_2880_420 0 0.008f
c2517 net8_M3_2880_500 0 0.008f
r1289 net8_M3_2880_500 net8_M3_2880_504 0.16
c2518 net8_M3_2880_500 0 0.0004f
c2519 net8_M3_2880_504 0 0.0004f
r1290 net8_M3_2880_504 net8_M3_2880_584 3.2
c2520 net8_M3_2880_504 0 0.008f
c2521 net8_M3_2880_584 0 0.008f
r1291 net8_M3_2880_584 net8_M3_2880_624 1.6
c2522 net8_M3_2880_584 0 0.004f
c2523 net8_M3_2880_624 0 0.004f
r1292 vss_M3_560_132 vss_M3_560_168 1.44
c2524 vss_M3_560_132 0 0.0036f
c2525 vss_M3_560_168 0 0.0036f
r1293 vss_M3_560_168 vss_M3_560_248 3.2
c2526 vss_M3_560_168 0 0.008f
c2527 vss_M3_560_248 0 0.008f
r1294 vss_M3_560_248 vss_M3_560_328 3.2
c2528 vss_M3_560_248 0 0.008f
c2529 vss_M3_560_328 0 0.008f
r1295 vss_M3_560_328 vss_M3_560_408 3.2
c2530 vss_M3_560_328 0 0.008f
c2531 vss_M3_560_408 0 0.008f
r1296 vss_M3_560_408 vss_M3_560_420 0.48
c2532 vss_M3_560_408 0 0.0012000000000000001f
c2533 vss_M3_560_420 0 0.0012000000000000001f
r1297 vss_M3_560_420 vss_M3_560_456 1.44
c2534 vss_M3_560_420 0 0.0036f
c2535 vss_M3_560_456 0 0.0036f
r1298 vss_M3_800_132 vss_M3_800_168 1.44
c2536 vss_M3_800_132 0 0.0036f
c2537 vss_M3_800_168 0 0.0036f
r1299 vss_M3_800_168 vss_M3_800_248 3.2
c2538 vss_M3_800_168 0 0.008f
c2539 vss_M3_800_248 0 0.008f
r1300 vss_M3_800_248 vss_M3_800_328 3.2
c2540 vss_M3_800_248 0 0.008f
c2541 vss_M3_800_328 0 0.008f
r1301 vss_M3_800_328 vss_M3_800_408 3.2
c2542 vss_M3_800_328 0 0.008f
c2543 vss_M3_800_408 0 0.008f
r1302 vss_M3_800_408 vss_M3_800_420 0.48
c2544 vss_M3_800_408 0 0.0012000000000000001f
c2545 vss_M3_800_420 0 0.0012000000000000001f
r1303 vss_M3_800_420 vss_M3_800_456 1.44
c2546 vss_M3_800_420 0 0.0036f
c2547 vss_M3_800_456 0 0.0036f
r1304 id_M3_640__36 id_M3_640_0 1.44
c2548 id_M3_640__36 0 0.0036f
c2549 id_M3_640_0 0 0.0036f
r1305 id_M3_640_0 id_M3_640_80 3.2
c2550 id_M3_640_0 0 0.008f
c2551 id_M3_640_80 0 0.008f
r1306 id_M3_640_80 id_M3_640_160 3.2
c2552 id_M3_640_80 0 0.008f
c2553 id_M3_640_160 0 0.008f
r1307 id_M3_640_160 id_M3_640_240 3.2
c2554 id_M3_640_160 0 0.008f
c2555 id_M3_640_240 0 0.008f
r1308 id_M3_640_240 id_M3_640_252 0.48
c2556 id_M3_640_240 0 0.0012000000000000001f
c2557 id_M3_640_252 0 0.0012000000000000001f
r1309 id_M3_640_252 id_M3_640_332 3.2
c2558 id_M3_640_252 0 0.008f
c2559 id_M3_640_332 0 0.008f
r1310 id_M3_640_332 id_M3_640_412 3.2
c2560 id_M3_640_332 0 0.008f
c2561 id_M3_640_412 0 0.008f
r1311 id_M3_640_412 id_M3_640_492 3.2
c2562 id_M3_640_412 0 0.008f
c2563 id_M3_640_492 0 0.008f
r1312 id_M3_640_492 id_M3_640_504 0.48
c2564 id_M3_640_492 0 0.0012000000000000001f
c2565 id_M3_640_504 0 0.0012000000000000001f
r1313 id_M3_640_504 id_M3_640_540 1.44
c2566 id_M3_640_504 0 0.0036f
c2567 id_M3_640_540 0 0.0036f
r1314 id_M3_880_216 id_M3_880_252 1.44
c2568 id_M3_880_216 0 0.0036f
c2569 id_M3_880_252 0 0.0036f
r1315 id_M3_880_252 id_M3_880_332 3.2
c2570 id_M3_880_252 0 0.008f
c2571 id_M3_880_332 0 0.008f
r1316 id_M3_880_332 id_M3_880_412 3.2
c2572 id_M3_880_332 0 0.008f
c2573 id_M3_880_412 0 0.008f
r1317 id_M3_880_412 id_M3_880_492 3.2
c2574 id_M3_880_412 0 0.008f
c2575 id_M3_880_492 0 0.008f
r1318 id_M3_880_492 id_M3_880_504 0.48
c2576 id_M3_880_492 0 0.0012000000000000001f
c2577 id_M3_880_504 0 0.0012000000000000001f
r1319 id_M3_880_504 id_M3_880_540 1.44
c2578 id_M3_880_504 0 0.0036f
c2579 id_M3_880_540 0 0.0036f
r1320 net10_M3_720_300 net10_M3_720_336 1.44
c2580 net10_M3_720_300 0 0.0036f
c2581 net10_M3_720_336 0 0.0036f
r1321 net10_M3_720_336 net10_M3_720_416 3.2
c2582 net10_M3_720_336 0 0.008f
c2583 net10_M3_720_416 0 0.008f
r1322 net10_M3_720_416 net10_M3_720_496 3.2
c2584 net10_M3_720_416 0 0.008f
c2585 net10_M3_720_496 0 0.008f
r1323 net10_M3_720_496 net10_M3_720_576 3.2
c2586 net10_M3_720_496 0 0.008f
c2587 net10_M3_720_576 0 0.008f
r1324 net10_M3_720_576 net10_M3_720_588 0.48
c2588 net10_M3_720_576 0 0.0012000000000000001f
c2589 net10_M3_720_588 0 0.0012000000000000001f
r1325 net10_M3_720_588 net10_M3_720_624 1.44
c2590 net10_M3_720_588 0 0.0036f
c2591 net10_M3_720_624 0 0.0036f
r1326 net10_M3_960_128 net10_M3_960_208 3.2
c2592 net10_M3_960_128 0 0.008f
c2593 net10_M3_960_208 0 0.008f
r1327 net10_M3_960_208 net10_M3_960_288 3.2
c2594 net10_M3_960_208 0 0.008f
c2595 net10_M3_960_288 0 0.008f
r1328 net10_M3_960_288 net10_M3_960_336 1.92
c2596 net10_M3_960_288 0 0.0048000000000000004f
c2597 net10_M3_960_336 0 0.0048000000000000004f
r1329 net10_M3_960_336 net10_M3_960_416 3.2
c2598 net10_M3_960_336 0 0.008f
c2599 net10_M3_960_416 0 0.008f
r1330 net10_M3_960_416 net10_M3_960_496 3.2
c2600 net10_M3_960_416 0 0.008f
c2601 net10_M3_960_496 0 0.008f
r1331 net10_M3_960_496 net10_M3_960_576 3.2
c2602 net10_M3_960_496 0 0.008f
c2603 net10_M3_960_576 0 0.008f
r1332 net10_M3_960_576 net10_M3_960_588 0.48
c2604 net10_M3_960_576 0 0.0012000000000000001f
c2605 net10_M3_960_588 0 0.0012000000000000001f
r1333 net10_M3_960_168 net10_M3_960_248 3.2
c2606 net10_M3_960_168 0 0.008f
c2607 net10_M3_960_248 0 0.008f
r1334 net10_M3_960_248 net10_M3_960_328 3.2
c2608 net10_M3_960_248 0 0.008f
c2609 net10_M3_960_328 0 0.008f
r1335 net10_M3_960_328 net10_M3_960_408 3.2
c2610 net10_M3_960_328 0 0.008f
c2611 net10_M3_960_408 0 0.008f
r1336 net10_M3_960_408 net10_M3_960_488 3.2
c2612 net10_M3_960_408 0 0.008f
c2613 net10_M3_960_488 0 0.008f
r1337 net10_M3_960_488 net10_M3_960_568 3.2
c2614 net10_M3_960_488 0 0.008f
c2615 net10_M3_960_568 0 0.008f
r1338 net10_M3_960_568 net10_M3_960_624 2.24
c2616 net10_M3_960_568 0 0.005600000000000001f
c2617 net10_M3_960_624 0 0.005600000000000001f
r1339 net8_M3_2160_216 net8_M3_2160_252 1.44
c2618 net8_M3_2160_216 0 0.0036f
c2619 net8_M3_2160_252 0 0.0036f
r1340 net8_M3_2160_252 net8_M3_2160_332 3.2
c2620 net8_M3_2160_252 0 0.008f
c2621 net8_M3_2160_332 0 0.008f
r1341 net8_M3_2160_332 net8_M3_2160_412 3.2
c2622 net8_M3_2160_332 0 0.008f
c2623 net8_M3_2160_412 0 0.008f
r1342 net8_M3_2160_412 net8_M3_2160_492 3.2
c2624 net8_M3_2160_412 0 0.008f
c2625 net8_M3_2160_492 0 0.008f
r1343 net8_M3_2160_492 net8_M3_2160_504 0.48
c2626 net8_M3_2160_492 0 0.0012000000000000001f
c2627 net8_M3_2160_504 0 0.0012000000000000001f
r1344 net8_M3_2160_504 net8_M3_2160_544 1.6
c2628 net8_M3_2160_504 0 0.004f
c2629 net8_M3_2160_544 0 0.004f
r1345 vdd_M3_3600_231 vdd_M3_3600_311 3.2
c2630 vdd_M3_3600_231 0 0.008f
c2631 vdd_M3_3600_311 0 0.008f
r1346 vdd_M3_3600_311 vdd_M3_3600_336 1.0
c2632 vdd_M3_3600_311 0 0.0025000000000000005f
c2633 vdd_M3_3600_336 0 0.0025000000000000005f
r1347 vdd_M3_3600_336 vdd_M3_3600_416 3.2
c2634 vdd_M3_3600_336 0 0.008f
c2635 vdd_M3_3600_416 0 0.008f
r1348 vdd_M3_3600_416 vdd_M3_3600_441 1.0
c2636 vdd_M3_3600_416 0 0.0025000000000000005f
c2637 vdd_M3_3600_441 0 0.0025000000000000005f
r1349 vdd_M3_3360_231 vdd_M3_3360_311 3.2
c2638 vdd_M3_3360_231 0 0.008f
c2639 vdd_M3_3360_311 0 0.008f
r1350 vdd_M3_3360_311 vdd_M3_3360_336 1.0
c2640 vdd_M3_3360_311 0 0.0025000000000000005f
c2641 vdd_M3_3360_336 0 0.0025000000000000005f
r1351 vdd_M3_3360_336 vdd_M3_3360_416 3.2
c2642 vdd_M3_3360_336 0 0.008f
c2643 vdd_M3_3360_416 0 0.008f
r1352 vdd_M3_3360_416 vdd_M3_3360_441 1.0
c2644 vdd_M3_3360_416 0 0.0025000000000000005f
c2645 vdd_M3_3360_441 0 0.0025000000000000005f
r1353 vout_M3_2480_48 vout_M3_2480_84 1.44
c2646 vout_M3_2480_48 0 0.0036f
c2647 vout_M3_2480_84 0 0.0036f
r1354 vout_M3_2480_84 vout_M3_2480_164 3.2
c2648 vout_M3_2480_84 0 0.008f
c2649 vout_M3_2480_164 0 0.008f
r1355 vout_M3_2480_164 vout_M3_2480_244 3.2
c2650 vout_M3_2480_164 0 0.008f
c2651 vout_M3_2480_244 0 0.008f
r1356 vout_M3_2480_244 vout_M3_2480_324 3.2
c2652 vout_M3_2480_244 0 0.008f
c2653 vout_M3_2480_324 0 0.008f
r1357 vout_M3_2480_324 vout_M3_2480_336 0.48
c2654 vout_M3_2480_324 0 0.0012000000000000001f
c2655 vout_M3_2480_336 0 0.0012000000000000001f
r1358 vout_M3_2480_252 vout_M3_2480_332 3.2
c2656 vout_M3_2480_252 0 0.008f
c2657 vout_M3_2480_332 0 0.008f
r1359 vout_M3_2480_332 vout_M3_2480_372 1.6
c2658 vout_M3_2480_332 0 0.004f
c2659 vout_M3_2480_372 0 0.004f
r1360 vout_M3_2640_147 vout_M3_2640_227 3.2
c2660 vout_M3_2640_147 0 0.008f
c2661 vout_M3_2640_227 0 0.008f
r1361 vout_M3_2640_227 vout_M3_2640_252 1.0
c2662 vout_M3_2640_227 0 0.0025000000000000005f
c2663 vout_M3_2640_252 0 0.0025000000000000005f
r1362 vout_M3_2640_252 vout_M3_2640_332 3.2
c2664 vout_M3_2640_252 0 0.008f
c2665 vout_M3_2640_332 0 0.008f
r1363 vout_M3_2640_332 vout_M3_2640_357 1.0
c2666 vout_M3_2640_332 0 0.0025000000000000005f
c2667 vout_M3_2640_357 0 0.0025000000000000005f
r1364 vout_M3_2400__36 vout_M3_2400_0 1.44
c2668 vout_M3_2400__36 0 0.0036f
c2669 vout_M3_2400_0 0 0.0036f
r1365 vout_M3_2400_0 vout_M3_2400_80 3.2
c2670 vout_M3_2400_0 0 0.008f
c2671 vout_M3_2400_80 0 0.008f
r1366 vout_M3_2400_80 vout_M3_2400_160 3.2
c2672 vout_M3_2400_80 0 0.008f
c2673 vout_M3_2400_160 0 0.008f
r1367 vout_M3_2400_160 vout_M3_2400_240 3.2
c2674 vout_M3_2400_160 0 0.008f
c2675 vout_M3_2400_240 0 0.008f
r1368 vout_M3_2400_240 vout_M3_2400_252 0.48
c2676 vout_M3_2400_240 0 0.0012000000000000001f
c2677 vout_M3_2400_252 0 0.0012000000000000001f
r1369 vout_M3_2400_252 vout_M3_2400_288 1.44
c2678 vout_M3_2400_252 0 0.0036f
c2679 vout_M3_2400_288 0 0.0036f
r1370 net10_M3_1280_63 net10_M3_1280_143 3.2
c2680 net10_M3_1280_63 0 0.008f
c2681 net10_M3_1280_143 0 0.008f
r1371 net10_M3_1280_143 net10_M3_1280_168 1.0
c2682 net10_M3_1280_143 0 0.0025000000000000005f
c2683 net10_M3_1280_168 0 0.0025000000000000005f
r1372 net10_M3_1280_168 net10_M3_1280_248 3.2
c2684 net10_M3_1280_168 0 0.008f
c2685 net10_M3_1280_248 0 0.008f
r1373 net10_M3_1280_248 net10_M3_1280_273 1.0
c2686 net10_M3_1280_248 0 0.0025000000000000005f
c2687 net10_M3_1280_273 0 0.0025000000000000005f
r1374 vinp_M3_1920_128 vinp_M3_1920_208 3.2
c2688 vinp_M3_1920_128 0 0.008f
c2689 vinp_M3_1920_208 0 0.008f
r1375 vinp_M3_1920_208 vinp_M3_1920_288 3.2
c2690 vinp_M3_1920_208 0 0.008f
c2691 vinp_M3_1920_288 0 0.008f
r1376 vinp_M3_1920_288 vinp_M3_1920_368 3.2
c2692 vinp_M3_1920_288 0 0.008f
c2693 vinp_M3_1920_368 0 0.008f
r1377 vinp_M3_1920_368 vinp_M3_1920_420 2.08
c2694 vinp_M3_1920_368 0 0.0052f
c2695 vinp_M3_1920_420 0 0.0052f
r1378 vinp_M3_1920_168 vinp_M3_1920_248 3.2
c2696 vinp_M3_1920_168 0 0.008f
c2697 vinp_M3_1920_248 0 0.008f
r1379 vinp_M3_1920_248 vinp_M3_1920_328 3.2
c2698 vinp_M3_1920_248 0 0.008f
c2699 vinp_M3_1920_328 0 0.008f
r1380 vinp_M3_1920_328 vinp_M3_1920_408 3.2
c2700 vinp_M3_1920_328 0 0.008f
c2701 vinp_M3_1920_408 0 0.008f
r1381 vinp_M3_1920_408 vinp_M3_1920_456 1.92
c2702 vinp_M3_1920_408 0 0.0048000000000000004f
c2703 vinp_M3_1920_456 0 0.0048000000000000004f
r1382 vinp_M3_1600__40 vinp_M3_1600_40 3.2
c2704 vinp_M3_1600__40 0 0.008f
c2705 vinp_M3_1600_40 0 0.008f
r1383 vinp_M3_1600_40 vinp_M3_1600_120 3.2
c2706 vinp_M3_1600_40 0 0.008f
c2707 vinp_M3_1600_120 0 0.008f
r1384 vinp_M3_1600_120 vinp_M3_1600_200 3.2
c2708 vinp_M3_1600_120 0 0.008f
c2709 vinp_M3_1600_200 0 0.008f
r1385 vinp_M3_1600_200 vinp_M3_1600_252 2.08
c2710 vinp_M3_1600_200 0 0.0052f
c2711 vinp_M3_1600_252 0 0.0052f
r1386 vinp_M3_1600_0 vinp_M3_1600_80 3.2
c2712 vinp_M3_1600_0 0 0.008f
c2713 vinp_M3_1600_80 0 0.008f
r1387 vinp_M3_1600_80 vinp_M3_1600_160 3.2
c2714 vinp_M3_1600_80 0 0.008f
c2715 vinp_M3_1600_160 0 0.008f
r1388 vinp_M3_1600_160 vinp_M3_1600_240 3.2
c2716 vinp_M3_1600_160 0 0.008f
c2717 vinp_M3_1600_240 0 0.008f
r1389 vinp_M3_1600_240 vinp_M3_1600_288 1.92
c2718 vinp_M3_1600_240 0 0.0048000000000000004f
c2719 vinp_M3_1600_288 0 0.0048000000000000004f
r1390 vinp_M3_1360__36 vinp_M3_1360_0 1.44
c2720 vinp_M3_1360__36 0 0.0036f
c2721 vinp_M3_1360_0 0 0.0036f
r1391 vinp_M3_1360_0 vinp_M3_1360_80 3.2
c2722 vinp_M3_1360_0 0 0.008f
c2723 vinp_M3_1360_80 0 0.008f
r1392 vinp_M3_1360_80 vinp_M3_1360_160 3.2
c2724 vinp_M3_1360_80 0 0.008f
c2725 vinp_M3_1360_160 0 0.008f
r1393 vinp_M3_1360_160 vinp_M3_1360_240 3.2
c2726 vinp_M3_1360_160 0 0.008f
c2727 vinp_M3_1360_240 0 0.008f
r1394 vinp_M3_1360_240 vinp_M3_1360_252 0.48
c2728 vinp_M3_1360_240 0 0.0012000000000000001f
c2729 vinp_M3_1360_252 0 0.0012000000000000001f
r1395 vinp_M3_1360_252 vinp_M3_1360_288 1.44
c2730 vinp_M3_1360_252 0 0.0036f
c2731 vinp_M3_1360_288 0 0.0036f
r1396 vdd_M2_3920_0 vdd_M3_3920_0 50
r1397 vdd_M2_3920_168 vdd_M3_3920_168 50
r1398 vdd_M2_3920_336 vdd_M3_3920_336 50
r1399 vdd_M2_3760_168 vdd_M3_3760_168 50
r1400 vdd_M2_3760_336 vdd_M3_3760_336 50
r1401 net8_M2_3840_252 net8_M3_3840_252 50
r1402 net8_M2_3840_420 net8_M3_3840_420 50
r1403 net8_M2_3680_252 net8_M3_3680_252 50
r1404 net8_M2_3680_420 net8_M3_3680_420 50
r1405 vdd_M2_3280_168 vdd_M3_3280_168 50
r1406 vdd_M2_3280_420 vdd_M3_3280_420 50
r1407 vdd_M2_3040_168 vdd_M3_3040_168 50
r1408 vdd_M2_3040_420 vdd_M3_3040_420 50
r1409 vout_M2_3200_252 vout_M3_3200_252 50
r1410 vout_M2_3200_504 vout_M3_3200_504 50
r1411 vout_M2_2960_84 vout_M3_2960_84 50
r1412 vout_M2_2960_252 vout_M3_2960_252 50
r1413 vout_M2_2960_504 vout_M3_2960_504 50
r1414 net8_M2_3120_336 net8_M3_3120_336 50
r1415 net8_M2_3120_588 net8_M3_3120_588 50
r1416 net8_M2_2880_336 net8_M3_2880_336 50
r1417 net8_M2_2880_588 net8_M3_2880_588 50
r1418 vss_M2_560_168 vss_M3_560_168 50
r1419 vss_M2_560_420 vss_M3_560_420 50
r1420 vss_M2_800_168 vss_M3_800_168 50
r1421 vss_M2_800_420 vss_M3_800_420 50
r1422 id_M2_640_0 id_M3_640_0 50
r1423 id_M2_640_252 id_M3_640_252 50
r1424 id_M2_640_504 id_M3_640_504 50
r1425 id_M2_880_252 id_M3_880_252 50
r1426 id_M2_880_504 id_M3_880_504 50
r1427 net10_M2_720_336 net10_M3_720_336 50
r1428 net10_M2_720_588 net10_M3_720_588 50
r1429 net10_M2_960_336 net10_M3_960_336 50
r1430 net10_M2_960_588 net10_M3_960_588 50
r1431 net8_M2_2160_252 net8_M3_2160_252 50
r1432 vdd_M2_3360_336 vdd_M3_3360_336 50
r1433 vdd_M2_3600_336 vdd_M3_3600_336 50
r1434 vout_M2_2400_0 vout_M3_2400_0 50
r1435 vout_M2_2400_252 vout_M3_2400_252 50
r1436 vout_M2_2480_84 vout_M3_2480_84 50
r1437 vout_M2_2480_336 vout_M3_2480_336 50
r1438 vout_M2_2640_252 vout_M3_2640_252 50
r1439 net10_M2_1280_168 net10_M3_1280_168 50
r1440 vinp_M2_1360_0 vinp_M3_1360_0 50
r1441 vinp_M2_1360_252 vinp_M3_1360_252 50
r1442 vinp_M2_1600_252 vinp_M3_1600_252 50
r1443 vinp_M2_1920_420 vinp_M3_1920_420 50
r1444 net8_M4_2840_420 net8_M4_2880_420 1.2
c2732 net8_M4_2840_420 0 0.004f
c2733 net8_M4_2880_420 0 0.004f
r1445 net8_M4_2880_420 net8_M4_2960_420 2.4
c2734 net8_M4_2880_420 0 0.008f
c2735 net8_M4_2960_420 0 0.008f
r1446 net8_M4_2960_420 net8_M4_3040_420 2.4
c2736 net8_M4_2960_420 0 0.008f
c2737 net8_M4_3040_420 0 0.008f
r1447 net8_M4_3040_420 net8_M4_3120_420 2.4
c2738 net8_M4_3040_420 0 0.008f
c2739 net8_M4_3120_420 0 0.008f
r1448 net8_M4_3120_420 net8_M4_3200_420 2.4
c2740 net8_M4_3120_420 0 0.008f
c2741 net8_M4_3200_420 0 0.008f
r1449 net8_M4_3200_420 net8_M4_3280_420 2.4
c2742 net8_M4_3200_420 0 0.008f
c2743 net8_M4_3280_420 0 0.008f
r1450 net8_M4_3280_420 net8_M4_3360_420 2.4
c2744 net8_M4_3280_420 0 0.008f
c2745 net8_M4_3360_420 0 0.008f
r1451 net8_M4_3360_420 net8_M4_3440_420 2.4
c2746 net8_M4_3360_420 0 0.008f
c2747 net8_M4_3440_420 0 0.008f
r1452 net8_M4_3440_420 net8_M4_3520_420 2.4
c2748 net8_M4_3440_420 0 0.008f
c2749 net8_M4_3520_420 0 0.008f
r1453 net8_M4_3520_420 net8_M4_3600_420 2.4
c2750 net8_M4_3520_420 0 0.008f
c2751 net8_M4_3600_420 0 0.008f
r1454 net8_M4_3600_420 net8_M4_3680_420 2.4
c2752 net8_M4_3600_420 0 0.008f
c2753 net8_M4_3680_420 0 0.008f
r1455 net8_M4_3680_420 net8_M4_3720_420 1.2
c2754 net8_M4_3680_420 0 0.004f
c2755 net8_M4_3720_420 0 0.004f
r1456 net8_M4_2120_504 net8_M4_2160_504 1.2
c2756 net8_M4_2120_504 0 0.004f
c2757 net8_M4_2160_504 0 0.004f
r1457 net8_M4_2160_504 net8_M4_2240_504 2.4
c2758 net8_M4_2160_504 0 0.008f
c2759 net8_M4_2240_504 0 0.008f
r1458 net8_M4_2240_504 net8_M4_2320_504 2.4
c2760 net8_M4_2240_504 0 0.008f
c2761 net8_M4_2320_504 0 0.008f
r1459 net8_M4_2320_504 net8_M4_2400_504 2.4
c2762 net8_M4_2320_504 0 0.008f
c2763 net8_M4_2400_504 0 0.008f
r1460 net8_M4_2400_504 net8_M4_2480_504 2.4
c2764 net8_M4_2400_504 0 0.008f
c2765 net8_M4_2480_504 0 0.008f
r1461 net8_M4_2480_504 net8_M4_2560_504 2.4
c2766 net8_M4_2480_504 0 0.008f
c2767 net8_M4_2560_504 0 0.008f
r1462 net8_M4_2560_504 net8_M4_2640_504 2.4
c2768 net8_M4_2560_504 0 0.008f
c2769 net8_M4_2640_504 0 0.008f
r1463 net8_M4_2640_504 net8_M4_2720_504 2.4
c2770 net8_M4_2640_504 0 0.008f
c2771 net8_M4_2720_504 0 0.008f
r1464 net8_M4_2720_504 net8_M4_2800_504 2.4
c2772 net8_M4_2720_504 0 0.008f
c2773 net8_M4_2800_504 0 0.008f
r1465 net8_M4_2800_504 net8_M4_2880_504 2.4
c2774 net8_M4_2800_504 0 0.008f
c2775 net8_M4_2880_504 0 0.008f
r1466 net8_M4_2880_504 net8_M4_2920_504 1.2
c2776 net8_M4_2880_504 0 0.004f
c2777 net8_M4_2920_504 0 0.004f
r1467 vdd_M4_3000_336 vdd_M4_3040_336 1.2
c2778 vdd_M4_3000_336 0 0.004f
c2779 vdd_M4_3040_336 0 0.004f
r1468 vdd_M4_3040_336 vdd_M4_3120_336 2.4
c2780 vdd_M4_3040_336 0 0.008f
c2781 vdd_M4_3120_336 0 0.008f
r1469 vdd_M4_3120_336 vdd_M4_3200_336 2.4
c2782 vdd_M4_3120_336 0 0.008f
c2783 vdd_M4_3200_336 0 0.008f
r1470 vdd_M4_3200_336 vdd_M4_3280_336 2.4
c2784 vdd_M4_3200_336 0 0.008f
c2785 vdd_M4_3280_336 0 0.008f
r1471 vdd_M4_3280_336 vdd_M4_3360_336 2.4
c2786 vdd_M4_3280_336 0 0.008f
c2787 vdd_M4_3360_336 0 0.008f
r1472 vdd_M4_3360_336 vdd_M4_3400_336 1.2
c2788 vdd_M4_3360_336 0 0.004f
c2789 vdd_M4_3400_336 0 0.004f
r1473 vdd_M4_3560_336 vdd_M4_3600_336 1.2
c2790 vdd_M4_3560_336 0 0.004f
c2791 vdd_M4_3600_336 0 0.004f
r1474 vdd_M4_3600_336 vdd_M4_3680_336 2.4
c2792 vdd_M4_3600_336 0 0.008f
c2793 vdd_M4_3680_336 0 0.008f
r1475 vdd_M4_3680_336 vdd_M4_3760_336 2.4
c2794 vdd_M4_3680_336 0 0.008f
c2795 vdd_M4_3760_336 0 0.008f
r1476 vdd_M4_3760_336 vdd_M4_3800_336 1.2
c2796 vdd_M4_3760_336 0 0.004f
c2797 vdd_M4_3800_336 0 0.004f
r1477 vout_M4_2440_252 vout_M4_2480_252 1.2
c2798 vout_M4_2440_252 0 0.004f
c2799 vout_M4_2480_252 0 0.004f
r1478 vout_M4_2480_252 vout_M4_2560_252 2.4
c2800 vout_M4_2480_252 0 0.008f
c2801 vout_M4_2560_252 0 0.008f
r1479 vout_M4_2560_252 vout_M4_2640_252 2.4
c2802 vout_M4_2560_252 0 0.008f
c2803 vout_M4_2640_252 0 0.008f
r1480 vout_M4_2640_252 vout_M4_2680_252 1.2
c2804 vout_M4_2640_252 0 0.004f
c2805 vout_M4_2680_252 0 0.004f
r1481 net10_M4_920_168 net10_M4_960_168 1.2
c2806 net10_M4_920_168 0 0.004f
c2807 net10_M4_960_168 0 0.004f
r1482 net10_M4_960_168 net10_M4_1040_168 2.4
c2808 net10_M4_960_168 0 0.008f
c2809 net10_M4_1040_168 0 0.008f
r1483 net10_M4_1040_168 net10_M4_1120_168 2.4
c2810 net10_M4_1040_168 0 0.008f
c2811 net10_M4_1120_168 0 0.008f
r1484 net10_M4_1120_168 net10_M4_1200_168 2.4
c2812 net10_M4_1120_168 0 0.008f
c2813 net10_M4_1200_168 0 0.008f
r1485 net10_M4_1200_168 net10_M4_1280_168 2.4
c2814 net10_M4_1200_168 0 0.008f
c2815 net10_M4_1280_168 0 0.008f
r1486 net10_M4_1280_168 net10_M4_1320_168 1.2
c2816 net10_M4_1280_168 0 0.004f
c2817 net10_M4_1320_168 0 0.004f
r1487 vinp_M4_1400_168 vinp_M4_1480_168 2.4
c2818 vinp_M4_1400_168 0 0.008f
c2819 vinp_M4_1480_168 0 0.008f
r1488 vinp_M4_1480_168 vinp_M4_1560_168 2.4
c2820 vinp_M4_1480_168 0 0.008f
c2821 vinp_M4_1560_168 0 0.008f
r1489 vinp_M4_1560_168 vinp_M4_1640_168 2.4
c2822 vinp_M4_1560_168 0 0.008f
c2823 vinp_M4_1640_168 0 0.008f
r1490 vinp_M4_1640_168 vinp_M4_1720_168 2.4
c2824 vinp_M4_1640_168 0 0.008f
c2825 vinp_M4_1720_168 0 0.008f
r1491 vinp_M4_1720_168 vinp_M4_1800_168 2.4
c2826 vinp_M4_1720_168 0 0.008f
c2827 vinp_M4_1800_168 0 0.008f
r1492 vinp_M4_1800_168 vinp_M4_1880_168 2.4
c2828 vinp_M4_1800_168 0 0.008f
c2829 vinp_M4_1880_168 0 0.008f
r1493 vinp_M4_1880_168 vinp_M4_1920_168 1.2
c2830 vinp_M4_1880_168 0 0.004f
c2831 vinp_M4_1920_168 0 0.004f
r1494 vinp_M4_1440_168 vinp_M4_1520_168 2.4
c2832 vinp_M4_1440_168 0 0.008f
c2833 vinp_M4_1520_168 0 0.008f
r1495 vinp_M4_1520_168 vinp_M4_1600_168 2.4
c2834 vinp_M4_1520_168 0 0.008f
c2835 vinp_M4_1600_168 0 0.008f
r1496 vinp_M4_1600_168 vinp_M4_1680_168 2.4
c2836 vinp_M4_1600_168 0 0.008f
c2837 vinp_M4_1680_168 0 0.008f
r1497 vinp_M4_1680_168 vinp_M4_1760_168 2.4
c2838 vinp_M4_1680_168 0 0.008f
c2839 vinp_M4_1760_168 0 0.008f
r1498 vinp_M4_1760_168 vinp_M4_1840_168 2.4
c2840 vinp_M4_1760_168 0 0.008f
c2841 vinp_M4_1840_168 0 0.008f
r1499 vinp_M4_1840_168 vinp_M4_1920_168 2.4
c2842 vinp_M4_1840_168 0 0.008f
c2843 vinp_M4_1920_168 0 0.008f
r1500 vinp_M4_1920_168 vinp_M4_1960_168 1.2
c2844 vinp_M4_1920_168 0 0.004f
c2845 vinp_M4_1960_168 0 0.004f
r1501 vinp_M4_1400_0 vinp_M4_1480_0 2.4
c2846 vinp_M4_1400_0 0 0.008f
c2847 vinp_M4_1480_0 0 0.008f
r1502 vinp_M4_1480_0 vinp_M4_1560_0 2.4
c2848 vinp_M4_1480_0 0 0.008f
c2849 vinp_M4_1560_0 0 0.008f
r1503 vinp_M4_1560_0 vinp_M4_1600_0 1.2
c2850 vinp_M4_1560_0 0 0.004f
c2851 vinp_M4_1600_0 0 0.004f
r1504 vinp_M4_1440_0 vinp_M4_1520_0 2.4
c2852 vinp_M4_1440_0 0 0.008f
c2853 vinp_M4_1520_0 0 0.008f
r1505 vinp_M4_1520_0 vinp_M4_1600_0 2.4
c2854 vinp_M4_1520_0 0 0.008f
c2855 vinp_M4_1600_0 0 0.008f
r1506 vinp_M4_1600_0 vinp_M4_1640_0 1.2
c2856 vinp_M4_1600_0 0 0.004f
c2857 vinp_M4_1640_0 0 0.004f
r1507 net8_M3_2160_504 net8_M4_2160_504 50
r1508 net8_M3_2880_420 net8_M4_2880_420 50
r1509 net8_M3_2880_504 net8_M4_2880_504 50
r1510 net8_M3_3680_420 net8_M4_3680_420 50
r1511 vdd_M3_3040_336 vdd_M4_3040_336 50
r1512 vdd_M3_3360_336 vdd_M4_3360_336 50
r1513 vdd_M3_3600_336 vdd_M4_3600_336 50
r1514 vdd_M3_3760_336 vdd_M4_3760_336 50
r1515 vout_M3_2480_252 vout_M4_2480_252 50
r1516 vout_M3_2640_252 vout_M4_2640_252 50
r1517 net10_M3_960_168 net10_M4_960_168 50
r1518 net10_M3_1280_168 net10_M4_1280_168 50
r1519 vinp_M3_1600_0 vinp_M4_1600_0 50
r1520 vinp_M3_1920_168 vinp_M4_1920_168 50
r1521 vinp_M5_1440__40 vinp_M5_1440_0 0.8
c2858 vinp_M5_1440__40 0 0.004f
c2859 vinp_M5_1440_0 0 0.004f
r1522 vinp_M5_1440_0 vinp_M5_1440_80 1.6
c2860 vinp_M5_1440_0 0 0.008f
c2861 vinp_M5_1440_80 0 0.008f
r1523 vinp_M5_1440_80 vinp_M5_1440_160 1.6
c2862 vinp_M5_1440_80 0 0.008f
c2863 vinp_M5_1440_160 0 0.008f
r1524 vinp_M5_1440_160 vinp_M5_1440_168 0.16
c2864 vinp_M5_1440_160 0 0.0008f
c2865 vinp_M5_1440_168 0 0.0008f
r1525 vinp_M5_1440_168 vinp_M5_1440_208 0.8
c2866 vinp_M5_1440_168 0 0.004f
c2867 vinp_M5_1440_208 0 0.004f
r1526 vinp_M4_1440_0 vinp_M5_1440_0 50
r1527 vinp_M4_1440_168 vinp_M5_1440_168 50
r1528 net_m1_M1_X0_Y0_G net8_M1_3840_168 50
r1529 net_m1_M1_X0_Y0_S vdd_M1_3920_336 50
r1530 net_m1_M1_X0_Y0_S vdd_M1_3920_462 50
r1531 net_m1_M1_X0_Y0_S vdd_M1_3920_588 50
r1532 net_m1_M1_X0_Y0_D net8_M1_3760_336 50
r1533 net_m1_M1_X0_Y0_D net8_M1_3760_462 50
r1534 net_m1_M1_X0_Y0_D net8_M1_3760_588 50
r1535 net_m2_M1_X0_Y0_G net8_M1_3120_168 50
r1536 net_m2_M1_X0_Y0_S vdd_M1_3200_336 50
r1537 net_m2_M1_X0_Y0_S vdd_M1_3200_462 50
r1538 net_m2_M1_X0_Y0_S vdd_M1_3200_588 50
r1539 net_m2_M1_X0_Y0_D vout_M1_3040_336 50
r1540 net_m2_M1_X0_Y0_D vout_M1_3040_462 50
r1541 net_m2_M1_X0_Y0_D vout_M1_3040_588 50
r1542 net_m5_m4_M1_X0_Y0_G id_M1_400_168 50
r1543 net_m5_m4_M1_X0_Y0_S vss_M1_320_336 50
r1544 net_m5_m4_M1_X0_Y0_S vss_M1_320_462 50
r1545 net_m5_m4_M1_X0_Y0_S vss_M1_320_588 50
r1546 net_m5_m4_M1_X0_Y0_D id_M1_480_336 50
r1547 net_m5_m4_M1_X0_Y0_D id_M1_480_462 50
r1548 net_m5_m4_M1_X0_Y0_D id_M1_480_588 50
r1549 net_m5_m4_M2_X1_Y0_G id_M1_1040_168 50
r1550 net_m5_m4_M2_X1_Y0_S vss_M1_960_336 50
r1551 net_m5_m4_M2_X1_Y0_S vss_M1_960_462 50
r1552 net_m5_m4_M2_X1_Y0_S vss_M1_960_588 50
r1553 net_m5_m4_M2_X1_Y0_D net10_M1_1120_336 50
r1554 net_m5_m4_M2_X1_Y0_D net10_M1_1120_462 50
r1555 net_m5_m4_M2_X1_Y0_D net10_M1_1120_588 50
r1556 net_m0_m3_M1_X0_Y0_G vinp_M1_1760_168 50
r1557 net_m0_m3_M1_X0_Y0_S net10_M1_1680_336 50
r1558 net_m0_m3_M1_X0_Y0_S net10_M1_1680_462 50
r1559 net_m0_m3_M1_X0_Y0_S net10_M1_1680_588 50
r1560 net_m0_m3_M1_X0_Y0_D net8_M1_1840_336 50
r1561 net_m0_m3_M1_X0_Y0_D net8_M1_1840_462 50
r1562 net_m0_m3_M1_X0_Y0_D net8_M1_1840_588 50
r1563 net_m0_m3_M2_X1_Y0_G vinn_M1_2400_168 50
r1564 net_m0_m3_M2_X1_Y0_S net10_M1_2320_336 50
r1565 net_m0_m3_M2_X1_Y0_S net10_M1_2320_462 50
r1566 net_m0_m3_M2_X1_Y0_S net10_M1_2320_588 50
r1567 net_m0_m3_M2_X1_Y0_D vout_M1_2480_336 50
r1568 net_m0_m3_M2_X1_Y0_D vout_M1_2480_462 50
r1569 net_m0_m3_M2_X1_Y0_D vout_M1_2480_588 50
x1_M1_X0_Y0_0 net_m1_M1_X0_Y0_D net_m1_M1_X0_Y0_G net_m1_M1_X0_Y0_diff vdd! PMOS l=2e-08 nfin=12 w=2.7e-07
x1_M1_X0_Y0_1 net_m1_M1_X0_Y0_diff net_m1_M1_X0_Y0_G net_m1_M1_X0_Y0_S vdd! PMOS l=2e-08 nfin=12 w=2.7e-07
x2_M1_X0_Y0_0 net_m2_M1_X0_Y0_D net_m2_M1_X0_Y0_G net_m2_M1_X0_Y0_diff vdd! PMOS l=2e-08 nfin=12 w=2.7e-07
x2_M1_X0_Y0_1 net_m2_M1_X0_Y0_diff net_m2_M1_X0_Y0_G net_m2_M1_X0_Y0_S vdd! PMOS l=2e-08 nfin=12 w=2.7e-07
x5_m4_M1_X0_Y0_0 net_m5_m4_M1_X0_Y0_D net_m5_m4_M1_X0_Y0_G net_m5_m4_M1_X0_Y0_diff gnd! NMOS l=2e-08 nfin=12 w=2.7e-07
x5_m4_M1_X0_Y0_1 net_m5_m4_M1_X0_Y0_diff net_m5_m4_M1_X0_Y0_G net_m5_m4_M1_X0_Y0_S gnd! NMOS l=2e-08 nfin=12 w=2.7e-07
x5_m4_M2_X1_Y0_0 net_m5_m4_M2_X1_Y0_D net_m5_m4_M2_X1_Y0_G net_m5_m4_M2_X1_Y0_diff gnd! NMOS l=2e-08 nfin=12 w=2.7e-07
x5_m4_M2_X1_Y0_1 net_m5_m4_M2_X1_Y0_diff net_m5_m4_M2_X1_Y0_G net_m5_m4_M2_X1_Y0_S gnd! NMOS l=2e-08 nfin=12 w=2.7e-07
x0_m3_M1_X0_Y0_0 net_m0_m3_M1_X0_Y0_D net_m0_m3_M1_X0_Y0_G net_m0_m3_M1_X0_Y0_diff gnd! NMOS l=2e-08 nfin=12 w=2.7e-07
x0_m3_M1_X0_Y0_1 net_m0_m3_M1_X0_Y0_diff net_m0_m3_M1_X0_Y0_G net_m0_m3_M1_X0_Y0_S gnd! NMOS l=2e-08 nfin=12 w=2.7e-07
x0_m3_M2_X1_Y0_0 net_m0_m3_M2_X1_Y0_D net_m0_m3_M2_X1_Y0_G net_m0_m3_M2_X1_Y0_diff gnd! NMOS l=2e-08 nfin=12 w=2.7e-07
x0_m3_M2_X1_Y0_1 net_m0_m3_M2_X1_Y0_diff net_m0_m3_M2_X1_Y0_G net_m0_m3_M2_X1_Y0_S gnd! NMOS l=2e-08 nfin=12 w=2.7e-07

**testbench
v2 vinp_M5_1440_0 0 DC 675e-3 AC 500e-3 180
v1 vinn_M2_2400_504 0 DC 675e-3 AC 500e-3
v0 vdd! 0 1000e-3
i5 vdd! id_M3_640_252 40e-6

cload vout_M4_2440_252 0 350e-15

.AC DEC 100 1.0 1e11

.PRINT AC vdb(vout_M4_2440_252)

.END
